.include /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical


.param  sw_stat_mismatch = 0
.param  sw_stat_global = 0

.include ../netlist/Programmable_2stage_opamp_wo_res_pex.spice
X1 vout vout_t vbiasp vbiasn vin2 vin1 vprog vss vdd opamp2

V1 vdd GND 3.3
V2 vss GND 0
V3 vin1 GND dc 0.8 ac 1
V4 vin2 GND dc 0.8 ac 0 
V5 vprog GND dc 0
V6 vbiasp GND dc 0.9
V7 vbiasn GND dc 1



.save i(v1)
.save i(v2)
.save i(v3)
.save i(v4)
.save i(v5)
.save all

.control

let begin = 1
let step = 0.1
let final = 1
let test = begin
let cnt = 0
let ind = ((final-begin)/step)
let n = vector(ind)
let power = vector(ind)

set color0 = white
set color1 = black
set hcopydevtype = svg
setcs svg_stropts = ( black Arial Arial )
set nolegend

set inoise = ' '


let test = begin
while test le final

    alter @v5[dc] = test
    print @v5[dc]
    let test = test + step

    op

    let ic = v1#branch
    let power[cnt] = 3.3*(-ic)
    print power[cnt]
    let cnt = cnt + 1

end




let test = begin
let cnt = 0
while test le final

    alter @v5[dc] = test
    print @v5[dc]
    let test = test + step

    noise v(vout) v3 dec 100 20K 2MEG 1

    let n[cnt] = inoise_total
    let cnt = cnt + 1
    setplot previous
    set inoise = ( $inoise ({$curplot}.inoise_spectrum) )

end



plot $inoise xlabel Frequency ylabel Integrated_Noise(uV) title Integrated_Noise
plot n vs power xlabel Power(mW) ylabel Integrated_Noise(uV) title 'OTA_2stage Integrated_Noise_vs_Power'

hardcopy ../output/Noise.svg $inoise xlabel  Frequency(Hz) ylabel Integrated_Noise(uV) title 'OTA_2stage Integrated_Noise'
hardcopy ../output/Noise_vs_Power.svg n vs power xlabel Power(mW) ylabel Integrated_Noise(uV) title 'OTA_2stage Integrated_Noise_vs_Power'

print n

.endc


.GLOBAL GND

.end

* NGSPICE file created from opamp2_nodw.ext - technology: gf180mcuC

.subckt opamp2 vout vout_t vbiasp vbiasn vin2 vin1 vprog vss vdd
X0 vss a_31806_2835# vout vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X1 a_13786_2835# vin2.t0 a_7580_3503# vdd.t556 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X2 vss vss.t226 vss vss nfet_03v3 ad=367.68p pd=0.00156024 as=2.6p ps=10.52u w=10u l=300n
X3 a_13786_2835# vin2.t1 a_7580_3503# vdd.t555 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X4 vout a_31806_2835# vss vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X5 a_13786_5007# vin1.t0 a_7580_3503# vdd.t521 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X6 a_19749_n2296# vin1.t1 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X7 vdd vdd.t364 vdd vdd.t155 pfet_03v3 ad=463.44p pd=0.0020616 as=1.1p ps=5.88u w=2.5u l=3u
X8 a_7580_3503# vin1.t2 a_13786_5007# vdd.t552 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X9 a_9856_n4071# vin1.t3 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X10 vdd vdd.t360 vdd vdd.t16 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X11 a_11312_n4152# a_6084_4175# a_6084_4175# vss nfet_03v3 ad=520f pd=2.52u as=880f ps=4.88u w=2u l=1000n
X12 vdd vdd.t356 vdd vdd.t331 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X13 a_13786_2835# a_31806_5067# vss vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=1000n
X14 a_9856_n4071# vin2.t2 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X15 a_7580_3503# a_5796_5519# vdd vdd.t21 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X16 vdd vdd.t351 vdd vdd.t352 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X17 a_7580_3503# vin2.t3 a_13786_2835# vdd.t554 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X18 a_19749_n6676# vin2.t4 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X19 vdd a_28902_5067# vout vdd.t326 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X20 a_19749_n6676# vin2.t5 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X21 a_9656_n5262# a_5010_6963# a_5010_6963# vss nfet_03v3 ad=520f pd=2.52u as=880f ps=4.88u w=2u l=1000n
X22 vout_t vdd.t601 vout vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X23 a_13786_5007# vin1.t4 a_7580_3503# vdd.t556 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X24 vdd vdd.t347 vdd vdd.t6 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X25 vss vss.t222 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X26 a_9856_n4071# vin2.t6 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X27 vout a_28902_5067# vdd vdd.t321 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X28 a_9656_n5262# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X29 a_7580_3503# vin2.t7 a_13786_2835# vdd.t553 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X30 vss vss.t218 vss vss nfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X31 a_7580_3503# vin2.t8 a_13786_2835# vdd.t552 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X32 vdd vdd.t343 vdd vdd.t115 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X33 vss vss.t214 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X34 vss a_31806_2835# vout vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X35 a_7580_3503# vin1.t5 a_13786_5007# vdd.t554 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X36 vss vss.t210 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X37 a_19749_n2296# vin1.t6 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X38 vss vss.t206 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X39 vdd vdd.t339 vdd vdd.t308 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X40 vout vss.t308 vout_t vdd.t518 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X41 vdd vdd.t335 vdd vdd.t1 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X42 vss vss.t202 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X43 vout_t vdd.t606 vout vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X44 a_7580_3503# vin1.t7 a_13786_5007# vdd.t553 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X45 a_19749_n6676# vin2.t9 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X46 a_5010_6963# a_5010_6963# a_9656_n5262# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X47 a_7580_3503# a_5796_5519# vdd vdd.t110 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X48 vdd vdd.t330 vdd vdd.t331 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X49 a_19749_n6676# vbiasp.t0 a_28902_5067# vdd.t558 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=3u
X50 vdd a_21261_4878# a_19749_n6676# vdd.t369 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X51 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X52 a_11312_n4152# a_11312_n4152# vss vss nfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=1000n
X53 vdd vdd.t325 vdd vdd.t326 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X54 a_13786_2835# vin2.t10 a_7580_3503# vdd.t551 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X55 a_9856_n4071# vin1.t8 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X56 a_13786_2835# vin2.t11 a_7580_3503# vdd.t550 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X57 vout vdd.t609 vout_t vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X58 a_19749_n6676# vin2.t12 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X59 a_7580_3503# a_5796_5519# vdd vdd.t97 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X60 a_7580_3503# a_5796_5519# vdd vdd.t1 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X61 a_7580_3503# vin1.t9 a_13786_5007# vdd.t549 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X62 vss vss.t198 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X63 vdd vdd.t320 vdd vdd.t321 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X64 a_19749_n2296# vin1.t10 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X65 a_5796_5519# a_5796_5519# vdd vdd.t494 pfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=3u
X66 vss a_31806_2835# vout vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X67 vdd vdd.t316 vdd vdd.t291 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X68 vdd a_28902_5067# vout vdd.t286 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X69 vdd a_21261_4878# a_19749_n2296# vdd.t410 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X70 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X71 vdd vdd.t312 vdd vdd.t155 pfet_03v3 ad=1.1p pd=5.88u as=0 ps=0 w=2.5u l=3u
X72 vdd a_28902_5067# vout vdd.t281 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X73 vss vss.t194 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X74 a_4788_4131# a_4788_4131# a_4700_4175# vdd.t137 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X75 a_13786_5007# vin1.t11 a_7580_3503# vdd.t548 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X76 a_13786_5007# vin1.t12 a_7580_3503# vdd.t551 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X77 a_7580_3503# a_5796_5519# vdd vdd.t1 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X78 a_9656_n5262# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=1000n
X79 vss vss.t190 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X80 a_13786_5007# vin1.t13 a_7580_3503# vdd.t550 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X81 vdd vdd.t307 vdd vdd.t308 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X82 a_19749_n6676# vin2.t13 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X83 a_9856_n4071# vin2.t14 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X84 vdd vdd.t303 vdd vdd.t115 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X85 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X86 vss vss.t186 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X87 a_7580_3503# vin2.t15 a_13786_2835# vdd.t549 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X88 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=1000n
X89 a_28902_5067# vout.t36 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X90 a_19749_n6676# vin2.t16 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X91 a_9856_n4071# vin2.t17 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X92 vdd vdd.t299 vdd vdd.t264 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X93 a_7580_3503# a_5796_5519# vdd vdd.t155 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X94 a_7580_3503# a_5796_5519# vdd vdd.t69 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X95 a_13786_2835# vin2.t18 a_7580_3503# vdd.t548 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X96 a_7580_3503# a_5796_5519# vdd vdd.t1 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X97 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X98 a_9856_n4071# vin2.t19 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X99 a_19749_n2296# vin1.t14 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X100 vdd vdd.t295 vdd vdd.t115 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X101 a_13786_5007# a_31806_5067# vss vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=1000n
X102 a_7580_3503# a_5796_5519# vdd vdd.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X103 vss vss.t182 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X104 vdd vprog.t0 a_5010_6963# vdd.t594 pfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=3u
X105 a_13786_5007# vin1.t15 a_7580_3503# vdd.t547 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X106 a_11512_n3371# a_5010_6963# a_4788_4131# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X107 vdd vdd.t290 vdd vdd.t291 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X108 vdd vdd.t285 vdd vdd.t286 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X109 vss vss.t178 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X110 a_9856_n4071# vin2.t20 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X111 a_19749_n6676# a_21261_4878# vdd vdd.t407 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X112 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X113 vdd vdd.t280 vdd vdd.t281 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X114 a_9856_n4071# vin1.t16 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X115 a_7580_3503# a_5796_5519# vdd vdd.t110 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X116 vout_t vss.t316 vout vdd.t517 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X117 vdd vdd.t276 vdd vdd.t115 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X118 vss vss.t174 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X119 vss vss.t170 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X120 a_31806_2835# a_4788_4131# a_28902_5067# vdd.t557 pfet_03v3 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=1000n
X121 vss vss.t166 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X122 vss vss.t162 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X123 a_28902_5067# vout.t35 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X124 a_6084_4175# a_6084_4175# a_11312_n4152# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X125 vdd vdd.t272 vdd vdd.t250 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X126 vdd a_28902_5067# vout vdd.t245 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X127 a_7580_3503# a_5796_5519# vdd vdd.t97 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X128 vdd a_21261_4878# a_19749_n6676# vdd.t410 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X129 a_4788_4131# a_4788_4131# a_4700_4175# vdd.t83 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X130 a_13786_2835# vin2.t21 a_7580_3503# vdd.t547 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X131 a_13786_5007# vin1.t17 a_7580_3503# vdd.t546 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X132 a_9856_n4071# vin1.t18 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X133 a_19749_n2296# vin1.t19 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X134 a_13786_5007# vin1.t20 a_7580_3503# vdd.t545 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X135 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=1000n
X136 a_7580_3503# a_5796_5519# vdd vdd.t110 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X137 vdd vdd.t268 vdd vdd.t115 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X138 vout_t vdd.t623 vout vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X139 vdd vdd.t263 vdd vdd.t264 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X140 a_9856_n4071# vin1.t21 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X141 vout_t vss.t321 vout vdd.t516 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X142 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=1000n
X143 vdd vdd.t259 vdd vdd.t240 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X144 a_19749_n2296# vin1.t22 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X145 a_7580_3503# a_5796_5519# vdd vdd.t21 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X146 a_7580_3503# a_5796_5519# vdd vdd.t97 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X147 a_9856_n4071# vin1.t23 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X148 vss vss.t158 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X149 a_19749_n6676# vin2.t22 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X150 a_13786_2835# vin2.t23 a_7580_3503# vdd.t546 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X151 vdd vdd.t254 vdd vdd.t255 pfet_03v3 ad=0 pd=0 as=880f ps=4.88u w=2u l=3u
X152 a_19749_n2296# vin1.t24 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X153 a_13786_2835# vin2.t24 a_7580_3503# vdd.t545 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X154 vout a_28902_5067# vdd vdd.t235 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X155 a_7580_3503# a_5796_5519# vdd vdd.t69 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X156 a_31806_2835# vbiasn.t0 a_13786_2835# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=1000n
X157 vout vss.t323 vout_t vdd.t515 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X158 a_7580_3503# vin2.t25 a_13786_2835# vdd.t544 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X159 a_5010_6963# a_5010_6963# a_9656_n5262# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X160 a_19749_n6676# vbiasp.t1 a_28902_5067# vdd.t368 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=3u
X161 a_7580_3503# vin1.t25 a_13786_5007# vdd.t543 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X162 vss vss.t154 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X163 a_5884_4131# a_5884_4131# a_5796_5519# vdd.t264 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X164 a_13786_5007# vin1.t26 a_7580_3503# vdd.t542 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X165 vss a_31806_2835# vout vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X166 vdd vdd.t249 vdd vdd.t250 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X167 vout_t vdd.t628 vout vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X168 a_7580_3503# a_5796_5519# vdd vdd.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X169 vdd vdd.t244 vdd vdd.t245 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X170 vout a_28902_5067# vdd vdd.t226 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X171 a_19749_n2296# a_21261_4878# vdd vdd.t407 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X172 a_9856_n4071# vin2.t26 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X173 a_19749_n6676# vin2.t27 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X174 a_5884_4131# a_5884_4131# a_5796_5519# vdd.t264 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X175 a_7580_3503# vin1.t27 a_13786_5007# vdd.t544 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X176 a_31806_5067# a_4788_4131# a_21261_4878# vdd.t557 pfet_03v3 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=1000n
X177 a_7580_3503# a_5796_5519# vdd vdd.t69 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X178 a_7580_3503# vin2.t28 a_13786_2835# vdd.t543 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X179 vout vdd.t630 vout_t vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X180 a_13786_2835# vin2.t29 a_7580_3503# vdd.t542 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X181 a_31806_2835# vout.t3 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X182 vss vss.t150 vss vss nfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X183 a_19749_n2296# a_21261_4878# vdd vdd.t400 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X184 a_21261_4878# vbiasp.t2 a_19749_n2296# vdd.t559 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X185 a_7580_3503# a_5796_5519# vdd vdd.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X186 a_9656_n5262# a_5010_6963# a_5010_6963# vss nfet_03v3 ad=880f pd=4.88u as=520f ps=2.52u w=2u l=1000n
X187 a_13786_5007# vin1.t28 a_7580_3503# vdd.t541 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X188 vout a_31806_2835# vss vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X189 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X190 vdd vdd.t239 vdd vdd.t240 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X191 vss vss.t146 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X192 a_6084_4175# a_5884_4131# a_5796_4175# vdd.t264 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X193 vdd vdd.t234 vdd vdd.t235 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X194 a_9856_n4071# vin1.t29 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X195 vss vss.t142 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X196 vout a_31806_2835# vss vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X197 a_11512_n3371# a_5010_6963# a_4788_4131# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X198 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=1000n
X199 vss vss.t138 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X200 vout vdd.t633 vout_t vss nfet_03v3 ad=260f pd=1.52u as=440f ps=2.88u w=1000n l=280n
X201 vdd vdd.t230 vdd vdd.t209 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X202 a_7580_3503# vin1.t30 a_13786_5007# vdd.t539 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X203 a_9856_n4071# vin1.t31 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X204 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=1000n
X205 a_7580_3503# a_5796_5519# vdd vdd.t21 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X206 a_13786_2835# vin2.t30 a_7580_3503# vdd.t541 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X207 vdd vdd.t225 vdd vdd.t226 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X208 a_7580_3503# vin2.t31 a_13786_2835# vdd.t540 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X209 vss a_9656_n5262# a_9656_n5262# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X210 a_6084_4175# a_6084_4175# a_11312_n4152# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X211 a_5884_4131# a_5884_4131# a_5796_5519# vdd.t240 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X212 a_19749_n2296# vbiasp.t3 a_21261_4878# vdd.t368 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=3u
X213 a_13786_5007# vin1.t32 a_7580_3503# vdd.t538 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X214 a_19749_n2296# vin1.t33 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X215 vdd vdd.t221 vdd vdd.t196 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X216 vout a_28902_5067# vdd vdd.t191 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X217 a_7580_3503# vin2.t32 a_13786_2835# vdd.t539 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X218 a_19749_n2296# vin1.t34 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X219 vdd a_21261_4878# a_19749_n6676# vdd.t397 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=3u
X220 a_28902_5067# vout.t34 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X221 a_5010_6963# a_5010_6963# a_9656_n5262# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X222 a_9856_n4071# vin1.t35 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X223 a_7580_3503# a_5796_5519# vdd vdd.t21 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X224 a_5884_4131# a_5884_4131# a_5796_5519# vdd.t240 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X225 a_7580_3503# vin1.t36 a_13786_5007# vdd.t535 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X226 a_9856_n4071# vin2.t33 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X227 a_7580_3503# a_5796_5519# vdd vdd.t1 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X228 a_7580_3503# vin1.t37 a_13786_5007# vdd.t540 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X229 vss vss.t134 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X230 vout_t vss.t330 vout vdd.t514 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X231 vss vss.t130 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X232 a_13786_2835# vin2.t34 a_7580_3503# vdd.t538 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X233 a_13786_2835# vin2.t35 a_7580_3503# vdd.t537 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X234 a_13786_2835# vin2.t36 a_7580_3503# vdd.t536 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X235 a_19749_n2296# vin1.t38 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X236 vdd vdd.t217 vdd vdd.t137 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X237 vss vss.t126 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X238 vout vdd.t638 vout_t vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X239 a_19749_n6676# a_21261_4878# vdd vdd.t400 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X240 a_11072_n909# a_9656_n5262# vss vss nfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=1000n
X241 vss vss.t122 vss vss nfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X242 a_28902_5067# vbiasp.t4 a_19749_n6676# vdd.t559 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X243 vdd vdd.t213 vdd vdd.t177 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X244 vdd vdd.t208 vdd vdd.t209 pfet_03v3 ad=2.6p pd=10.52u as=0 ps=0 w=10u l=300n
X245 a_31806_5067# vbiasn.t1 a_13786_5007# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=1000n
X246 a_9856_n4071# vin2.t37 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X247 a_19749_n6676# vin2.t38 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X248 vdd vdd.t204 vdd vdd.t172 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X249 a_7580_3503# vin2.t39 a_13786_2835# vdd.t535 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X250 a_6084_4175# a_5884_4131# a_5796_4175# vdd.t240 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X251 vout_t vdd.t642 vout vss nfet_03v3 ad=440f pd=2.88u as=260f ps=1.52u w=1000n l=280n
X252 a_13786_5007# vin1.t39 a_7580_3503# vdd.t537 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X253 a_13786_5007# vin1.t40 a_7580_3503# vdd.t536 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X254 vdd vdd.t200 vdd vdd.t155 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X255 vout_t vss.t334 vout vdd.t513 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X256 a_19749_n6676# vin2.t40 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X257 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=1000n
X258 vdd vdd.t195 vdd vdd.t196 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X259 a_9856_n4071# vin2.t41 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X260 a_9856_n4071# vin1.t41 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X261 a_7580_3503# vin2.t42 a_13786_2835# vdd.t505 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X262 a_19749_n2296# vin1.t42 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X263 vdd vdd.t190 vdd vdd.t191 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X264 a_19749_n6676# vin2.t43 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X265 a_7580_3503# vin2.t44 a_13786_2835# vdd.t534 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X266 vss a_31806_5067# a_13786_2835# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=1000n
X267 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X268 vdd vdd.t185 vdd vdd.t186 pfet_03v3 ad=0 pd=0 as=880f ps=4.88u w=2u l=3u
X269 vout vss.t335 vout_t vdd.t512 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X270 a_31806_2835# vout.t2 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X271 vdd vdd.t181 vdd vdd.t142 pfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X272 vss vss.t118 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X273 a_19749_n6676# vin2.t45 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X274 vss vss.t114 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X275 a_19749_n6676# vin2.t46 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X276 a_9656_n5262# a_5010_6963# a_5010_6963# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X277 a_7580_3503# vin2.t47 a_13786_2835# vdd.t533 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X278 vout_t vdd.t648 vout vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X279 a_7580_3503# vin1.t43 a_13786_5007# vdd.t505 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X280 vdd a_21261_4878# a_19749_n2296# vdd.t397 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=3u
X281 vss a_9656_n5262# a_9656_n5262# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X282 a_7580_3503# vin1.t44 a_13786_5007# vdd.t506 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X283 a_7580_3503# vin1.t45 a_13786_5007# vdd.t534 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X284 vdd vdd.t176 vdd vdd.t177 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X285 vdd vdd.t171 vdd vdd.t172 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X286 a_19749_n2296# vin1.t46 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X287 vdd vdd.t167 vdd vdd.t137 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X288 a_7580_3503# a_5796_5519# vdd vdd.t1 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X289 a_11072_n909# a_5010_6963# a_5884_4131# vss nfet_03v3 ad=151.6f pd=1.64u as=151.6f ps=1.64u w=220n l=1000n
X290 a_9856_n4071# vin1.t47 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X291 vdd vdd.t163 vdd vdd.t83 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X292 vout vss.t338 vout_t vdd.t511 pfet_03v3 ad=520f pd=2.52u as=880f ps=4.88u w=2u l=280n
X293 vdd a_21261_4878# a_19749_n6676# vdd.t392 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X294 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X295 a_7580_3503# vin1.t48 a_13786_5007# vdd.t533 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X296 vdd vdd.t159 vdd vdd.t110 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X297 vdd a_28902_5067# vout vdd.t120 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X298 a_7580_3503# vin2.t48 a_13786_2835# vdd.t506 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X299 vss vss.t110 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X300 a_9856_n4071# vin2.t49 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X301 vss vss.t106 vss vss nfet_03v3 ad=0 pd=0 as=2.2p ps=10.88u w=5u l=1000n
X302 vdd vdd.t154 vdd vdd.t155 pfet_03v3 ad=1.1p pd=5.88u as=0 ps=0 w=2.5u l=3u
X303 a_13786_2835# vin2.t50 a_7580_3503# vdd.t532 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X304 vdd vdd.t150 vdd vdd.t137 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X305 a_7580_3503# a_5796_5519# vdd vdd.t1 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X306 a_13786_5007# vin1.t49 a_7580_3503# vdd.t531 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X307 vdd vdd.t146 vdd vdd.t97 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X308 a_5796_4175# a_5796_5519# vdd vdd.t453 pfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=3u
X309 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X310 vss vss.t102 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X311 a_9856_n4071# vin2.t51 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X312 vdd vdd.t141 vdd vdd.t142 pfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X313 vss vss.t98 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X314 vdd vdd.t136 vdd vdd.t137 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X315 a_9856_n4071# vin1.t50 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X316 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X317 a_7580_3503# a_5796_5519# vdd vdd.t155 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X318 a_13786_5007# vin1.t51 a_7580_3503# vdd.t532 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X319 a_13786_2835# vin2.t52 a_7580_3503# vdd.t531 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X320 a_9656_n5262# a_5010_6963# a_5010_6963# vss nfet_03v3 ad=520f pd=2.52u as=880f ps=4.88u w=2u l=1000n
X321 a_9856_n4071# vin2.t53 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X322 vss vss.t94 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X323 vout a_28902_5067# vdd vdd.t88 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X324 a_19749_n6676# vin2.t54 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X325 vout vss.t344 vout_t vdd.t510 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X326 a_7580_3503# vin2.t55 a_13786_2835# vdd.t530 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X327 a_31806_5067# a_6084_4175# a_21261_4878# vss nfet_03v3 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=1000n
X328 a_4788_4131# a_5010_6963# a_11512_n3371# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X329 a_19749_n6676# vin2.t56 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X330 a_9856_n4071# vin2.t57 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X331 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X332 a_9856_n4071# vin1.t52 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X333 vdd vdd.t132 vdd vdd.t69 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X334 a_7580_3503# a_5796_5519# vdd vdd.t155 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X335 vdd vdd.t128 vdd vdd.t78 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X336 vdd vdd.t124 vdd vdd.t83 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X337 vdd vdd.t119 vdd vdd.t120 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X338 a_4788_4131# a_4788_4131# a_4700_4175# vdd.t137 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X339 a_11312_n4152# a_6084_4175# a_6084_4175# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X340 vout_t vss.t345 vout vdd.t509 pfet_03v3 ad=880f pd=4.88u as=520f ps=2.52u w=2u l=280n
X341 vdd vdd.t114 vdd vdd.t115 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X342 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=1000n
X343 vdd vdd.t109 vdd vdd.t110 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X344 vdd vdd.t105 vdd vdd.t50 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X345 a_19749_n6676# vin2.t58 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X346 vdd a_4700_4175# a_4700_4175# vdd.t561 pfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=3u
X347 vss vss.t90 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X348 vdd vdd.t101 vdd vdd.t64 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X349 a_7580_3503# vin1.t53 a_13786_5007# vdd.t530 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X350 vdd a_21261_4878# a_19749_n2296# vdd.t392 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X351 vss vss.t86 vss vss nfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X352 vss a_31806_2835# vout vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X353 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=1000n
X354 vout vdd.t667 vout_t vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X355 vdd a_28902_5067# vout vdd.t55 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X356 a_19749_n6676# a_21261_4878# vdd vdd.t383 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X357 vss a_31806_5067# a_13786_5007# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=1000n
X358 a_13786_2835# vin2.t59 a_7580_3503# vdd.t529 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X359 a_9656_n5262# a_5010_6963# a_5010_6963# vss nfet_03v3 ad=880f pd=4.88u as=520f ps=2.52u w=2u l=1000n
X360 vdd vdd.t96 vdd vdd.t97 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X361 a_19749_n2296# vin1.t54 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X362 a_7580_3503# a_5796_5519# vdd vdd.t155 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X363 vss vss.t82 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X364 vdd vdd.t92 vdd vdd.t83 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X365 vss vss.t78 vss vss nfet_03v3 ad=0 pd=0 as=1.76p ps=8.88u w=4u l=1000n
X366 a_4788_4131# a_5010_6963# a_11512_n3371# vss nfet_03v3 ad=880f pd=4.88u as=520f ps=2.52u w=2u l=1000n
X367 a_19749_n2296# a_21261_4878# vdd vdd.t378 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X368 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X369 a_7580_3503# vin2.t60 a_13786_2835# vdd.t528 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X370 a_9856_n4071# vin2.t61 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X371 vss vss.t74 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X372 vss vss.t70 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X373 a_7580_3503# a_5796_5519# vdd vdd.t110 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X374 vdd a_28902_5067# vout vdd.t45 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X375 vdd vdd.t87 vdd vdd.t88 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X376 vout_t vss.t352 vout vdd.t508 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X377 vdd a_28902_5067# vout vdd.t40 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X378 a_9856_n4071# vin2.t62 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X379 a_19749_n6676# vin2.t63 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X380 vdd vdd.t82 vdd vdd.t83 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=1000n
X381 a_11312_n4152# a_6084_4175# a_6084_4175# vss nfet_03v3 ad=880f pd=4.88u as=520f ps=2.52u w=2u l=1000n
X382 a_13786_5007# vin1.t55 a_7580_3503# vdd.t529 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X383 a_9856_n4071# vin2.t64 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X384 a_28902_5067# vout.t33 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X385 a_7580_3503# a_5796_5519# vdd vdd.t97 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X386 a_13786_2835# vbiasn.t2 a_31806_2835# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=1000n
X387 a_9856_n4071# vin1.t56 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X388 vdd vdd.t77 vdd vdd.t78 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X389 a_19749_n2296# vin1.t57 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X390 a_7580_3503# a_5796_5519# vdd vdd.t110 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X391 a_7580_3503# vin1.t58 a_13786_5007# vdd.t528 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X392 a_19749_n2296# vin1.t59 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X393 vdd vdd.t73 vdd vdd.t21 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X394 vdd vdd.t68 vdd vdd.t69 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X395 a_19749_n2296# vin1.t60 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X396 a_31806_2835# vout.t1 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X397 vss vss.t66 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X398 vout a_31806_2835# vss vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X399 a_7580_3503# a_5796_5519# vdd vdd.t97 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X400 vdd vdd.t63 vdd vdd.t64 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X401 vss vss.t62 vss vss nfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X402 vdd vdd.t59 vdd vdd.t31 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X403 a_28902_5067# vbiasp.t5 a_19749_n6676# vdd.t560 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=3u
X404 a_4788_4131# a_4788_4131# a_4700_4175# vdd.t83 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X405 vdd vdd.t54 vdd vdd.t55 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X406 vout a_28902_5067# vdd vdd.t26 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X407 vss vss.t58 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X408 vdd vdd.t49 vdd vdd.t50 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X409 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X410 vss vss.t54 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X411 a_6084_4175# a_5884_4131# a_5796_4175# vdd.t264 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X412 a_9856_n4071# vin2.t65 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X413 a_19749_n6676# vin2.t66 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X414 vss vss.t50 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X415 vdd a_21261_4878# a_19749_n6676# vdd.t375 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X416 a_7580_3503# a_5796_5519# vdd vdd.t110 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X417 a_7580_3503# vin1.t61 a_13786_5007# vdd.t525 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X418 a_7580_3503# a_5796_5519# vdd vdd.t69 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X419 a_13786_2835# vin2.t67 a_7580_3503# vdd.t527 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X420 vdd vdd.t44 vdd vdd.t45 pfet_03v3 ad=0 pd=0 as=4.4p ps=20.88u w=10u l=300n
X421 a_19749_n2296# a_21261_4878# vdd vdd.t383 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X422 vdd vdd.t39 vdd vdd.t40 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X423 a_7580_3503# a_5796_5519# vdd vdd.t97 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X424 a_9656_n5262# a_9656_n5262# vss vss nfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=1000n
X425 a_13786_2835# vin2.t68 a_7580_3503# vdd.t526 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X426 a_19749_n2296# a_21261_4878# vdd vdd.t372 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X427 a_19749_n2296# vin1.t62 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X428 a_9856_n4071# vin1.t63 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X429 a_7580_3503# a_5796_5519# vdd vdd.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X430 vdd vdd.t35 vdd vdd.t11 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X431 a_19749_n6676# a_21261_4878# vdd vdd.t378 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X432 a_7580_3503# vin1.t64 a_13786_5007# vdd.t523 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X433 a_7580_3503# a_5796_5519# vdd vdd.t69 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X434 a_9856_n4071# vin1.t65 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X435 vout vdd.t682 vout_t vss nfet_03v3 ad=260f pd=1.52u as=260f ps=1.52u w=1000n l=280n
X436 a_7580_3503# vin2.t69 a_13786_2835# vdd.t525 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X437 a_13786_5007# vin1.t66 a_7580_3503# vdd.t527 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X438 a_19749_n2296# vin1.t67 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X439 vss vss.t46 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X440 a_7580_3503# a_5796_5519# vdd vdd.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X441 a_19749_n6676# vin2.t70 a_9856_n4071# vss nfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X442 a_13786_5007# vin1.t68 a_7580_3503# vdd.t526 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X443 a_7580_3503# vin1.t69 a_13786_5007# vdd.t522 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X444 vdd vdd.t30 vdd vdd.t31 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X445 a_9856_n4071# vin2.t71 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X446 vss vss.t42 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X447 vdd vdd.t25 vdd vdd.t26 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X448 vdd vdd.t20 vdd vdd.t21 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X449 a_7580_3503# vin2.t72 a_13786_2835# vdd.t524 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X450 a_7580_3503# vin2.t73 a_13786_2835# vdd.t523 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=300n
X451 vss vss.t38 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X452 a_9856_n4071# vin1.t70 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=300n
X453 a_7580_3503# a_5796_5519# vdd vdd.t69 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X454 a_31806_2835# a_6084_4175# a_28902_5067# vss nfet_03v3 ad=4.4p pd=20.88u as=4.4p ps=20.88u w=10u l=1000n
X455 vout vss.t361 vout_t vdd.t507 pfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=280n
X456 a_13786_5007# vin1.t71 a_7580_3503# vdd.t520 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X457 a_19749_n2296# vin1.t72 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X458 a_9656_n5262# a_5010_6963# a_5010_6963# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X459 vdd vdd.t15 vdd vdd.t16 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X460 a_9856_n4071# vin1.t73 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X461 a_9856_n4071# vin2.t74 a_19749_n6676# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X462 vout a_28902_5067# vdd vdd.t352 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X463 a_21261_4878# vbiasp.t6 a_19749_n2296# vdd.t560 pfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=3u
X464 a_7580_3503# vin2.t75 a_13786_2835# vdd.t522 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X465 a_7580_3503# a_5796_5519# vdd vdd.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X466 a_19749_n2296# vin1.t74 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X467 a_6084_4175# a_5884_4131# a_5796_4175# vdd.t240 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=1000n
X468 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
X469 a_7580_3503# vin1.t75 a_13786_5007# vdd.t524 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X470 a_7580_3503# a_5796_5519# vdd vdd.t21 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X471 a_7580_3503# vin1.t76 a_13786_5007# vdd.t519 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X472 vdd vdd.t10 vdd vdd.t11 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X473 vdd a_21261_4878# a_19749_n2296# vdd.t375 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X474 a_31806_2835# vout.t0 cap_mim_2f0_m4m5_noshield c_width=25u c_length=25u
X475 a_5010_6963# a_5010_6963# a_9656_n5262# vss nfet_03v3 ad=520f pd=2.52u as=520f ps=2.52u w=2u l=1000n
X476 vdd vdd.t5 vdd vdd.t6 pfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X477 a_13786_5007# vin1.t77 a_7580_3503# vdd.t555 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X478 a_13786_2835# vin2.t76 a_7580_3503# vdd.t521 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X479 a_9856_n4071# vin1.t78 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X480 a_13786_2835# vin2.t77 a_7580_3503# vdd.t520 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X481 vss vss.t34 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X482 a_19749_n6676# vin2.t78 a_9856_n4071# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X483 a_13786_5007# vbiasn.t3 a_31806_5067# vss nfet_03v3 ad=2.6p pd=10.52u as=4.4p ps=20.88u w=10u l=1000n
X484 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=1000n
X485 a_11512_n3371# a_9656_n5262# vss vss nfet_03v3 ad=880f pd=4.88u as=880f ps=4.88u w=2u l=1000n
X486 a_9856_n4071# a_9656_n5262# vss vss nfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=1000n
X487 vss vss.t30 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X488 vdd vdd.t0 vdd vdd.t1 pfet_03v3 ad=0 pd=0 as=1.1p ps=5.88u w=2.5u l=3u
X489 a_7580_3503# a_5796_5519# vdd vdd.t21 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=3u
X490 a_19749_n6676# a_21261_4878# vdd vdd.t372 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X491 vss vss.t26 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X492 vout a_31806_2835# vss vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X493 vdd a_21261_4878# a_19749_n2296# vdd.t369 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=3u
X494 a_19749_n2296# vbiasp.t7 a_21261_4878# vdd.t558 pfet_03v3 ad=4.4p pd=20.88u as=2.6p ps=10.52u w=10u l=3u
X495 a_4788_4131# a_5010_6963# a_11512_n3371# vss nfet_03v3 ad=520f pd=2.52u as=880f ps=4.88u w=2u l=1000n
X496 a_7580_3503# vin2.t79 a_13786_2835# vdd.t519 pfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X497 a_9856_n4071# vin1.t79 a_19749_n2296# vss nfet_03v3 ad=2.6p pd=10.52u as=2.6p ps=10.52u w=10u l=300n
X498 vss vss.t22 vss vss nfet_03v3 ad=0 pd=0 as=2.6p ps=10.52u w=10u l=300n
X499 vss a_9656_n5262# a_9856_n4071# vss nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=1000n
R0 vout.n13 vout.n12 37.184
R1 vout.n15 vout.n14 12.737
R2 vout.n29 vout.n28 5.457
R3 vout.n10 pmos_3p3_CDNS_679510442370_0.S 3.513
R4 vout.n7 pmos_3p3_CDNS_679510442370_0.S 3.304
R5 vout.n10 pmos_3p3_CDNS_679510442370_0.S 3.135
R6 vout.n12 pmos_3p3_CDNS_679510442370_0.S 3.134
R7 vout.n9 pmos_3p3_CDNS_679510442370_0.S 3.134
R8 vout.n7 pmos_3p3_CDNS_679510442370_0.S 2.917
R9 vout.n11 pmos_3p3_CDNS_679510442370_0.S 2.914
R10 vout.n8 pmos_3p3_CDNS_679510442370_0.S 2.912
R11 vout.n14 vout 2.657
R12 vout.n27 vout.n23 2.361
R13 vout.n13 vout.n6 2.25
R14 vout.n0 vout 1.102
R15 vout.n18 nmos_3p3_CDNS_679510442372_0.S 0.911
R16 vout.n28 vout.n27 0.898
R17 vout.n19 vout.n18 0.626
R18 vout.n21 vout.n20 0.626
R19 vout.n22 vout.n21 0.626
R20 vout.n1 vout.n0 0.626
R21 vout.n31 vout.n30 0.626
R22 vout.n30 vout.n29 0.626
R23 vout.n14 vout.n13 0.5
R24 vout.n2 vout.t36 0.499
R25 vout.n29 vout 0.476
R26 vout.n30 vout 0.476
R27 vout.n31 vout 0.476
R28 vout.n1 vout 0.476
R29 vout.n0 vout 0.476
R30 vout.n6 vout.t2 0.446
R31 vout.n6 vout.t35 0.429
R32 vout.n23 vout.n22 0.41
R33 vout.n11 vout.n10 0.378
R34 vout.n8 vout.n7 0.378
R35 vout.n9 vout.n8 0.378
R36 vout.n12 vout.n9 0.378
R37 vout.n12 vout.n11 0.378
R38 nmos_3p3_CDNS_679510442372_0.S vout.n19 0.313
R39 vout.n20 nmos_3p3_CDNS_679510442372_0.S 0.313
R40 vout vout.n1 0.313
R41 vout vout.n31 0.313
R42 vout.n22 nmos_3p3_CDNS_679510442372_0.S 0.285
R43 vout.n21 nmos_3p3_CDNS_679510442372_0.S 0.285
R44 vout.n20 nmos_3p3_CDNS_679510442372_0.S 0.285
R45 vout.n19 nmos_3p3_CDNS_679510442372_0.S 0.285
R46 vout.n18 nmos_3p3_CDNS_679510442372_0.S 0.285
R47 vout.n4 vout.n3 0.116
R48 vout.t35 vout.n2 0.089
R49 vout.n3 vout.t1 0.069
R50 vout.t2 vout.n4 0.069
R51 vout.n3 vout.t0 0.065
R52 vout.n26 vout.n25 0.063
R53 vout.n17 vout.n16 0.063
R54 vout.n5 vout.t3 0.049
R55 vout.t2 vout.n5 0.039
R56 vout.n16 vout.n15 0.029
R57 vout.n28 vout.n17 0.029
R58 vout.n27 vout.n26 0.024
R59 vout.n25 vout.n24 0.024
R60 vout.t36 vout.t33 0.02
R61 vout.t33 vout.t34 0.019
R62 vss.n73 vss.t166 151.863
R63 vss.n77 vss.t150 151.863
R64 vss.n37 vss.t194 151.863
R65 vss.n41 vss.t218 151.863
R66 vss.n32 vss.t62 151.863
R67 vss.n57 vss.t206 151.863
R68 vss.n61 vss.t86 151.863
R69 vss.n52 vss.t122 151.863
R70 vss.n28 vss.t42 151.81
R71 vss.n48 vss.t50 151.81
R72 vss.n73 vss.t174 135.901
R73 vss.n74 vss.t102 135.901
R74 vss.n75 vss.t158 135.901
R75 vss.n76 vss.t222 135.901
R76 vss.n80 vss.t118 135.901
R77 vss.n79 vss.t178 135.901
R78 vss.n78 vss.t34 135.901
R79 vss.n77 vss.t110 135.901
R80 vss.n37 vss.t38 135.901
R81 vss.n38 vss.t154 135.901
R82 vss.n39 vss.t210 135.901
R83 vss.n40 vss.t90 135.901
R84 vss.n44 vss.t134 135.901
R85 vss.n43 vss.t198 135.901
R86 vss.n42 vss.t98 135.901
R87 vss.n41 vss.t146 135.901
R88 vss.n28 vss.t94 135.901
R89 vss.n29 vss.t202 135.901
R90 vss.n30 vss.t54 135.901
R91 vss.n31 vss.t126 135.901
R92 vss.n35 vss.t170 135.901
R93 vss.n34 vss.t46 135.901
R94 vss.n33 vss.t138 135.901
R95 vss.n32 vss.t190 135.901
R96 vss.n57 vss.t130 135.901
R97 vss.n58 vss.t226 135.901
R98 vss.n59 vss.t22 135.901
R99 vss.n60 vss.t142 135.901
R100 vss.n64 vss.t214 135.901
R101 vss.n63 vss.t66 135.901
R102 vss.n62 vss.t182 135.901
R103 vss.n61 vss.t26 135.901
R104 vss.n48 vss.t162 135.901
R105 vss.n49 vss.t70 135.901
R106 vss.n50 vss.t74 135.901
R107 vss.n51 vss.t186 135.901
R108 vss.n55 vss.t58 135.901
R109 vss.n54 vss.t114 135.901
R110 vss.n53 vss.t30 135.901
R111 vss.n52 vss.t82 135.901
R112 vss.n262 vss.t345 58.587
R113 vss.n267 vss.t338 58.587
R114 vss.n262 vss.t361 42.365
R115 vss.n263 vss.t330 42.365
R116 vss.n264 vss.t344 42.365
R117 vss.n265 vss.t316 42.365
R118 vss.n266 vss.t335 42.365
R119 vss.n271 vss.t352 42.365
R120 vss.n270 vss.t323 42.365
R121 vss.n269 vss.t334 42.365
R122 vss.n268 vss.t308 42.365
R123 vss.n267 vss.t321 42.365
R124 vss.n47 vss.t106 32.638
R125 vss.n47 vss.t78 22.87
R126 vss.n263 vss.n262 16.222
R127 vss.n264 vss.n263 16.222
R128 vss.n265 vss.n264 16.222
R129 vss.n266 vss.n265 16.222
R130 vss.n271 vss.n270 16.222
R131 vss.n270 vss.n269 16.222
R132 vss.n269 vss.n268 16.222
R133 vss.n268 vss.n267 16.222
R134 vss.n74 vss.n73 15.962
R135 vss.n75 vss.n74 15.962
R136 vss.n76 vss.n75 15.962
R137 vss.n80 vss.n79 15.962
R138 vss.n79 vss.n78 15.962
R139 vss.n78 vss.n77 15.962
R140 vss.n38 vss.n37 15.962
R141 vss.n39 vss.n38 15.962
R142 vss.n40 vss.n39 15.962
R143 vss.n44 vss.n43 15.962
R144 vss.n43 vss.n42 15.962
R145 vss.n42 vss.n41 15.962
R146 vss.n29 vss.n28 15.962
R147 vss.n30 vss.n29 15.962
R148 vss.n31 vss.n30 15.962
R149 vss.n35 vss.n34 15.962
R150 vss.n34 vss.n33 15.962
R151 vss.n33 vss.n32 15.962
R152 vss.n58 vss.n57 15.962
R153 vss.n59 vss.n58 15.962
R154 vss.n60 vss.n59 15.962
R155 vss.n64 vss.n63 15.962
R156 vss.n63 vss.n62 15.962
R157 vss.n62 vss.n61 15.962
R158 vss.n49 vss.n48 15.962
R159 vss.n50 vss.n49 15.962
R160 vss.n51 vss.n50 15.962
R161 vss.n55 vss.n54 15.962
R162 vss.n54 vss.n53 15.962
R163 vss.n53 vss.n52 15.962
R164 vss vss.n261 11.069
R165 vss.n81 vss.n80 8.662
R166 vss.n45 vss.n44 8.662
R167 vss.n65 vss.n64 8.662
R168 vss.n272 vss.n266 8.111
R169 vss.n272 vss.n271 8.111
R170 vss.n36 vss.n35 8.078
R171 vss.n56 vss.n55 8.078
R172 vss.n36 vss.n31 7.884
R173 vss.n56 vss.n51 7.884
R174 vss.n81 vss.n76 7.3
R175 vss.n45 vss.n40 7.3
R176 vss.n65 vss.n60 7.3
R177 vss.n67 vss.n66 6.119
R178 vss.n46 vss.n36 6.065
R179 vss.n66 vss.n56 6.065
R180 vss.n69 vss.n68 5.849
R181 vss.n261 vss.n260 5.844
R182 vss.n82 vss.n81 4.034
R183 vss.n46 vss.n45 4
R184 vss.n66 vss.n65 4
R185 vss vss.n272 4
R186 vss.n68 vss.n67 3.151
R187 vss.n258 vss.n257 2.868
R188 vss.n98 vss.n89 2.858
R189 vss.n145 vss.n105 2.555
R190 vss.n166 vss.n72 2.25
R191 vss.n187 vss.n71 2.25
R192 vss.n217 vss.n70 2.25
R193 vss.n227 vss.n69 2.25
R194 vss vss.n247 1.716
R195 vss.n146 vss.n82 1.401
R196 vss.n68 vss.n46 1.232
R197 vss.n259 vss.n258 1.121
R198 vss.n98 vss.n97 1.121
R199 vss.n98 vss.n93 1.121
R200 vss.n257 vss.n256 1.121
R201 vss.n105 vss.n104 1.121
R202 vss.n20 vss.n19 1.12
R203 vss.n88 vss.n8 1.12
R204 vss.n67 vss.n47 0.928
R205 vss.n201 vss.n200 0.563
R206 vss.n199 vss.n198 0.563
R207 vss.n197 vss.n196 0.563
R208 vss.n195 vss.n194 0.563
R209 vss.n187 vss.n186 0.563
R210 vss.n189 vss.n188 0.563
R211 vss.n191 vss.n190 0.563
R212 vss.n193 vss.n192 0.563
R213 vss.n203 vss.n202 0.563
R214 vss.n205 vss.n204 0.563
R215 vss.n207 vss.n206 0.563
R216 vss.n261 vss.n8 0.407
R217 vss.n248 vss 0.312
R218 vss.n247 vss.n246 0.087
R219 vss.n146 vss.n145 0.084
R220 vss.n145 vss.n144 0.062
R221 vss.n247 vss.n227 0.04
R222 vss.n139 vss.n138 0.02
R223 vss.n144 vss.n143 0.019
R224 vss.n143 vss.n142 0.019
R225 vss.n142 vss.n141 0.019
R226 vss.n141 vss.n140 0.019
R227 vss.n140 vss.n139 0.019
R228 vss.n138 vss.n137 0.019
R229 vss.n137 vss.n136 0.019
R230 vss.n136 vss.n135 0.019
R231 vss.n135 vss.n134 0.019
R232 vss.n134 vss.n133 0.019
R233 vss.n133 vss.n132 0.019
R234 vss.n132 vss.n131 0.019
R235 vss.n131 vss.n130 0.019
R236 vss.n130 vss.n129 0.019
R237 vss.n129 vss.n128 0.019
R238 vss.n128 vss.n127 0.019
R239 vss.n127 vss.n126 0.019
R240 vss.n126 vss.n125 0.019
R241 vss.n125 vss.n124 0.019
R242 vss.n124 vss.n123 0.019
R243 vss.n123 vss.n122 0.019
R244 vss.n122 vss.n121 0.019
R245 vss.n121 vss.n120 0.019
R246 vss.n120 vss.n119 0.019
R247 vss.n119 vss.n118 0.019
R248 vss.n118 vss.n117 0.019
R249 vss.n117 vss.n116 0.019
R250 vss.n116 vss.n115 0.019
R251 vss.n115 vss.n114 0.019
R252 vss.n114 vss.n113 0.019
R253 vss.n113 vss.n112 0.019
R254 vss.n112 vss.n111 0.019
R255 vss.n111 vss.n110 0.019
R256 vss.n110 vss.n109 0.019
R257 vss.n109 vss.n108 0.019
R258 vss.n108 vss.n107 0.019
R259 vss.n107 vss.n106 0.019
R260 vss.n229 vss.n228 0.019
R261 vss.n230 vss.n229 0.019
R262 vss.n231 vss.n230 0.019
R263 vss.n232 vss.n231 0.019
R264 vss.n233 vss.n232 0.019
R265 vss.n234 vss.n233 0.019
R266 vss.n235 vss.n234 0.019
R267 vss.n236 vss.n235 0.019
R268 vss.n237 vss.n236 0.019
R269 vss.n238 vss.n237 0.019
R270 vss.n239 vss.n238 0.019
R271 vss.n240 vss.n239 0.019
R272 vss.n241 vss.n240 0.019
R273 vss.n242 vss.n241 0.019
R274 vss.n243 vss.n242 0.019
R275 vss.n244 vss.n243 0.019
R276 vss.n245 vss.n244 0.019
R277 vss.n246 vss.n245 0.019
R278 vss.n86 vss.n85 0.016
R279 vss.n26 vss.n25 0.016
R280 vss.n17 vss.n16 0.014
R281 vss.n14 vss.n13 0.013
R282 vss.n7 vss.n6 0.013
R283 vss.n251 vss.n250 0.013
R284 vss.n258 vss.n21 0.013
R285 vss.n19 vss.n15 0.013
R286 vss.n103 vss.n102 0.013
R287 vss.n101 vss.n100 0.013
R288 vss.n24 vss.n23 0.013
R289 vss.n19 vss.n18 0.012
R290 vss.n100 vss.n99 0.012
R291 vss.n102 vss.n101 0.012
R292 vss.n23 vss.n22 0.012
R293 vss.n89 vss.n88 0.012
R294 vss.n88 vss.n87 0.012
R295 vss.n84 vss.n83 0.011
R296 vss.n104 vss.n98 0.011
R297 vss.n85 vss.n84 0.011
R298 vss.n104 vss.n103 0.011
R299 vss.n96 vss.n95 0.011
R300 vss.n249 vss.n248 0.011
R301 vss.n27 vss.n26 0.01
R302 vss.n257 vss.n27 0.01
R303 vss.n250 vss.n249 0.01
R304 vss.n2 vss.n1 0.01
R305 vss.n3 vss.n2 0.01
R306 vss.n6 vss.n5 0.01
R307 vss.n259 vss.n20 0.01
R308 vss.n12 vss.n11 0.01
R309 vss.n11 vss.n10 0.01
R310 vss.n260 vss.n259 0.01
R311 vss.n13 vss.n12 0.01
R312 vss.n10 vss.n9 0.01
R313 vss.n5 vss.n4 0.01
R314 vss.n1 vss.n0 0.01
R315 vss.n4 vss.n3 0.01
R316 vss.n93 vss.n90 0.01
R317 vss.n92 vss.n91 0.01
R318 vss.n97 vss.n94 0.01
R319 vss.n254 vss.n253 0.01
R320 vss.n256 vss.n254 0.01
R321 vss.n97 vss.n96 0.01
R322 vss.n93 vss.n92 0.01
R323 vss.n253 vss.n252 0.01
R324 vss.n256 vss.n255 0.01
R325 vss.n25 vss.n24 0.008
R326 vss.n87 vss.n86 0.008
R327 vss.n18 vss.n17 0.007
R328 vss.n8 vss.n7 0.007
R329 vss.n20 vss.n14 0.007
R330 vss.n252 vss.n251 0.007
R331 vss.n147 vss.n146 0.004
R332 vss.n148 vss.n147 0.004
R333 vss.n149 vss.n148 0.004
R334 vss.n150 vss.n149 0.004
R335 vss.n151 vss.n150 0.004
R336 vss.n152 vss.n151 0.004
R337 vss.n153 vss.n152 0.004
R338 vss.n154 vss.n153 0.004
R339 vss.n155 vss.n154 0.004
R340 vss.n156 vss.n155 0.004
R341 vss.n157 vss.n156 0.004
R342 vss.n158 vss.n157 0.004
R343 vss.n159 vss.n158 0.004
R344 vss.n160 vss.n159 0.004
R345 vss.n161 vss.n160 0.004
R346 vss.n162 vss.n161 0.004
R347 vss.n163 vss.n162 0.004
R348 vss.n164 vss.n163 0.004
R349 vss.n165 vss.n164 0.004
R350 vss.n167 vss.n166 0.004
R351 vss.n168 vss.n167 0.004
R352 vss.n169 vss.n168 0.004
R353 vss.n170 vss.n169 0.004
R354 vss.n171 vss.n170 0.004
R355 vss.n172 vss.n171 0.004
R356 vss.n173 vss.n172 0.004
R357 vss.n174 vss.n173 0.004
R358 vss.n175 vss.n174 0.004
R359 vss.n176 vss.n175 0.004
R360 vss.n177 vss.n176 0.004
R361 vss.n178 vss.n177 0.004
R362 vss.n179 vss.n178 0.004
R363 vss.n180 vss.n179 0.004
R364 vss.n181 vss.n180 0.004
R365 vss.n182 vss.n181 0.004
R366 vss.n183 vss.n182 0.004
R367 vss.n184 vss.n183 0.004
R368 vss.n185 vss.n184 0.004
R369 vss.n189 vss.n187 0.004
R370 vss.n191 vss.n189 0.004
R371 vss.n193 vss.n191 0.004
R372 vss.n195 vss.n193 0.004
R373 vss.n197 vss.n195 0.004
R374 vss.n199 vss.n197 0.004
R375 vss.n201 vss.n199 0.004
R376 vss.n203 vss.n201 0.004
R377 vss.n205 vss.n203 0.004
R378 vss.n207 vss.n205 0.004
R379 vss.n208 vss.n207 0.004
R380 vss.n209 vss.n208 0.004
R381 vss.n210 vss.n209 0.004
R382 vss.n211 vss.n210 0.004
R383 vss.n212 vss.n211 0.004
R384 vss.n213 vss.n212 0.004
R385 vss.n214 vss.n213 0.004
R386 vss.n215 vss.n214 0.004
R387 vss.n216 vss.n215 0.004
R388 vss.n218 vss.n217 0.004
R389 vss.n219 vss.n218 0.004
R390 vss.n220 vss.n219 0.004
R391 vss.n221 vss.n220 0.004
R392 vss.n222 vss.n221 0.004
R393 vss.n223 vss.n222 0.004
R394 vss.n224 vss.n223 0.004
R395 vss.n225 vss.n224 0.004
R396 vss.n226 vss.n225 0.004
R397 vss.n227 vss.n226 0.004
R398 vss.n166 vss.n165 0.003
R399 vss.n187 vss.n185 0.003
R400 vss.n217 vss.n216 0.003
R401 vin2.n29 vin2.n28 247.889
R402 vin2.n84 vin2.n38 212.639
R403 vin2.n19 vin2.t21 170.979
R404 vin2.n38 vin2.t69 158.774
R405 vin2.n37 vin2.t18 158.774
R406 vin2.n36 vin2.t79 158.774
R407 vin2.n35 vin2.t23 158.774
R408 vin2.n34 vin2.t28 158.774
R409 vin2.n33 vin2.t30 158.774
R410 vin2.n32 vin2.t39 158.774
R411 vin2.n31 vin2.t24 158.774
R412 vin2.n30 vin2.t48 158.774
R413 vin2.n29 vin2.t52 158.774
R414 vin2.n27 vin2.t73 158.774
R415 vin2.n26 vin2.t77 158.774
R416 vin2.n25 vin2.t75 158.774
R417 vin2.n24 vin2.t1 158.774
R418 vin2.n23 vin2.t8 158.774
R419 vin2.n22 vin2.t29 158.774
R420 vin2.n21 vin2.t15 158.774
R421 vin2.n20 vin2.t34 158.774
R422 vin2.n19 vin2.t32 158.774
R423 vin2.n39 vin2.t4 151.863
R424 vin2.n60 vin2.t70 151.863
R425 vin2.n48 vin2.t2 151.741
R426 vin2.n15 vin2.t10 144.743
R427 vin2.n0 vin2.t25 144.743
R428 vin2.n39 vin2.t62 135.901
R429 vin2.n40 vin2.t16 135.901
R430 vin2.n41 vin2.t65 135.901
R431 vin2.n42 vin2.t56 135.901
R432 vin2.n43 vin2.t26 135.901
R433 vin2.n44 vin2.t9 135.901
R434 vin2.n45 vin2.t37 135.901
R435 vin2.n46 vin2.t13 135.901
R436 vin2.n47 vin2.t71 135.901
R437 vin2.n60 vin2.t51 135.901
R438 vin2.n61 vin2.t22 135.901
R439 vin2.n62 vin2.t6 135.901
R440 vin2.n63 vin2.t45 135.901
R441 vin2.n64 vin2.t20 135.901
R442 vin2.n65 vin2.t78 135.901
R443 vin2.n66 vin2.t49 135.901
R444 vin2.n67 vin2.t5 135.901
R445 vin2.n68 vin2.t64 135.901
R446 vin2.n73 vin2.t63 135.901
R447 vin2.n74 vin2.t17 135.901
R448 vin2.n75 vin2.t66 135.901
R449 vin2.n76 vin2.t57 135.901
R450 vin2.n77 vin2.t27 135.901
R451 vin2.n78 vin2.t61 135.901
R452 vin2.n79 vin2.t38 135.901
R453 vin2.n80 vin2.t14 135.901
R454 vin2.n81 vin2.t46 135.901
R455 vin2.n82 vin2.t53 135.901
R456 vin2.n56 vin2.t43 135.779
R457 vin2.n55 vin2.t19 135.779
R458 vin2.n54 vin2.t58 135.779
R459 vin2.n53 vin2.t33 135.779
R460 vin2.n52 vin2.t12 135.779
R461 vin2.n51 vin2.t41 135.779
R462 vin2.n50 vin2.t40 135.779
R463 vin2.n49 vin2.t74 135.779
R464 vin2.n48 vin2.t54 135.779
R465 vin2.n15 vin2.t7 132.007
R466 vin2.n16 vin2.t59 132.007
R467 vin2.n17 vin2.t3 132.007
R468 vin2.n14 vin2.t76 132.007
R469 vin2.n13 vin2.t72 132.007
R470 vin2.n12 vin2.t67 132.007
R471 vin2.n11 vin2.t42 132.007
R472 vin2.n10 vin2.t35 132.007
R473 vin2.n9 vin2.t60 132.007
R474 vin2.n8 vin2.t0 132.007
R475 vin2.n7 vin2.t55 132.007
R476 vin2.n6 vin2.t50 132.007
R477 vin2.n5 vin2.t47 132.007
R478 vin2.n4 vin2.t68 132.007
R479 vin2.n3 vin2.t44 132.007
R480 vin2.n2 vin2.t36 132.007
R481 vin2.n1 vin2.t31 132.007
R482 vin2.n0 vin2.t11 132.007
R483 vin2.n28 vin2.n27 76.417
R484 vin2.n57 vin2.n47 54.937
R485 vin2.n83 vin2.n82 43.179
R486 vin2.n69 vin2.n68 43.176
R487 vin2.n73 vin2.n72 34.073
R488 vin2.n57 vin2.n56 33.956
R489 vin2.n9 vin2.n8 31.685
R490 vin2.n40 vin2.n39 15.962
R491 vin2.n41 vin2.n40 15.962
R492 vin2.n42 vin2.n41 15.962
R493 vin2.n43 vin2.n42 15.962
R494 vin2.n44 vin2.n43 15.962
R495 vin2.n45 vin2.n44 15.962
R496 vin2.n46 vin2.n45 15.962
R497 vin2.n47 vin2.n46 15.962
R498 vin2.n56 vin2.n55 15.962
R499 vin2.n55 vin2.n54 15.962
R500 vin2.n54 vin2.n53 15.962
R501 vin2.n53 vin2.n52 15.962
R502 vin2.n52 vin2.n51 15.962
R503 vin2.n51 vin2.n50 15.962
R504 vin2.n50 vin2.n49 15.962
R505 vin2.n49 vin2.n48 15.962
R506 vin2.n61 vin2.n60 15.962
R507 vin2.n62 vin2.n61 15.962
R508 vin2.n63 vin2.n62 15.962
R509 vin2.n64 vin2.n63 15.962
R510 vin2.n65 vin2.n64 15.962
R511 vin2.n66 vin2.n65 15.962
R512 vin2.n67 vin2.n66 15.962
R513 vin2.n68 vin2.n67 15.962
R514 vin2.n74 vin2.n73 15.962
R515 vin2.n75 vin2.n74 15.962
R516 vin2.n76 vin2.n75 15.962
R517 vin2.n77 vin2.n76 15.962
R518 vin2.n78 vin2.n77 15.962
R519 vin2.n79 vin2.n78 15.962
R520 vin2.n80 vin2.n79 15.962
R521 vin2.n81 vin2.n80 15.962
R522 vin2.n82 vin2.n81 15.962
R523 vin2 vin2.n84 15.653
R524 vin2.n28 vin2.n18 12.992
R525 vin2.n1 vin2.n0 12.736
R526 vin2.n2 vin2.n1 12.736
R527 vin2.n3 vin2.n2 12.736
R528 vin2.n4 vin2.n3 12.736
R529 vin2.n5 vin2.n4 12.736
R530 vin2.n6 vin2.n5 12.736
R531 vin2.n7 vin2.n6 12.736
R532 vin2.n8 vin2.n7 12.736
R533 vin2.n10 vin2.n9 12.736
R534 vin2.n11 vin2.n10 12.736
R535 vin2.n12 vin2.n11 12.736
R536 vin2.n13 vin2.n12 12.736
R537 vin2.n14 vin2.n13 12.736
R538 vin2.n17 vin2.n16 12.736
R539 vin2.n16 vin2.n15 12.736
R540 vin2.n38 vin2.n37 12.736
R541 vin2.n37 vin2.n36 12.736
R542 vin2.n36 vin2.n35 12.736
R543 vin2.n35 vin2.n34 12.736
R544 vin2.n34 vin2.n33 12.736
R545 vin2.n33 vin2.n32 12.736
R546 vin2.n32 vin2.n31 12.736
R547 vin2.n31 vin2.n30 12.736
R548 vin2.n30 vin2.n29 12.736
R549 vin2.n27 vin2.n26 12.736
R550 vin2.n26 vin2.n25 12.736
R551 vin2.n25 vin2.n24 12.736
R552 vin2.n24 vin2.n23 12.736
R553 vin2.n23 vin2.n22 12.736
R554 vin2.n22 vin2.n21 12.736
R555 vin2.n21 vin2.n20 12.736
R556 vin2.n20 vin2.n19 12.736
R557 vin2.n83 vin2.n57 11.152
R558 vin2.n18 vin2.n17 6.523
R559 vin2.n18 vin2.n14 6.212
R560 vin2.n84 vin2.n83 4.378
R561 vin2.n72 vin2.n71 1.492
R562 vin2.n70 vin2.n69 0.897
R563 vin2.n71 vin2.n59 0.027
R564 vin2.n72 vin2.n58 0.013
R565 vin2.n71 vin2.n70 0.009
R566 vdd.t110 vdd.t69 165.416
R567 vdd.t69 vdd.t50 165.416
R568 vdd.t97 vdd.t21 165.416
R569 vdd.t1 vdd.t97 165.416
R570 vdd.t558 vdd.t560 163.532
R571 vdd.n72 vdd.t44 146.95
R572 vdd.n67 vdd.t119 146.95
R573 vdd.n147 vdd.t181 146.95
R574 vdd.n138 vdd.t230 146.95
R575 vdd.n103 vdd.t141 146.95
R576 vdd.n94 vdd.t208 146.95
R577 vdd.n587 vdd.n583 140.833
R578 vdd.n72 vdd.t190 129.696
R579 vdd.n73 vdd.t280 129.696
R580 vdd.n74 vdd.t225 129.696
R581 vdd.n75 vdd.t325 129.696
R582 vdd.n76 vdd.t234 129.696
R583 vdd.n77 vdd.t244 129.696
R584 vdd.n78 vdd.t351 129.696
R585 vdd.n79 vdd.t285 129.696
R586 vdd.n67 vdd.t87 129.696
R587 vdd.n68 vdd.t54 129.696
R588 vdd.n69 vdd.t320 129.696
R589 vdd.n70 vdd.t39 129.696
R590 vdd.n147 vdd.t213 129.696
R591 vdd.n148 vdd.t221 129.696
R592 vdd.n149 vdd.t316 129.696
R593 vdd.n150 vdd.t339 129.696
R594 vdd.n138 vdd.t101 129.696
R595 vdd.n139 vdd.t128 129.696
R596 vdd.n140 vdd.t204 129.696
R597 vdd.n141 vdd.t59 129.696
R598 vdd.n142 vdd.t35 129.696
R599 vdd.n143 vdd.t15 129.696
R600 vdd.n144 vdd.t272 129.696
R601 vdd.n145 vdd.t5 129.696
R602 vdd.n103 vdd.t176 129.696
R603 vdd.n104 vdd.t195 129.696
R604 vdd.n105 vdd.t290 129.696
R605 vdd.n106 vdd.t307 129.696
R606 vdd.n94 vdd.t63 129.696
R607 vdd.n95 vdd.t77 129.696
R608 vdd.n96 vdd.t171 129.696
R609 vdd.n97 vdd.t30 129.696
R610 vdd.n98 vdd.t10 129.696
R611 vdd.n99 vdd.t360 129.696
R612 vdd.n100 vdd.t249 129.696
R613 vdd.n101 vdd.t347 129.696
R614 vdd.t368 vdd.t557 129.032
R615 vdd.n71 vdd.t25 127.621
R616 vdd.n102 vdd.t330 127.073
R617 vdd.n146 vdd.t356 127.066
R618 vdd.t560 vdd.t368 121.442
R619 vdd.t559 vdd.t558 121.442
R620 vdd.t378 vdd.t559 121.442
R621 vdd.t410 vdd.t378 121.442
R622 vdd.t372 vdd.t410 121.442
R623 vdd.t369 vdd.t372 121.442
R624 vdd.t400 vdd.t369 121.442
R625 vdd.n406 vdd.t525 99.706
R626 vdd.n377 vdd.t154 93.097
R627 vdd.n364 vdd.t200 92.205
R628 vdd.n378 vdd.n377 90.056
R629 vdd.n379 vdd.n378 90.056
R630 vdd.n380 vdd.n379 90.056
R631 vdd.n381 vdd.n380 90.056
R632 vdd.n382 vdd.n381 90.056
R633 vdd.n365 vdd.n364 89.164
R634 vdd.n366 vdd.n365 89.164
R635 vdd.n367 vdd.n366 89.164
R636 vdd.n368 vdd.n367 89.164
R637 vdd.n369 vdd.n368 89.164
R638 vdd.t83 vdd.t561 86.546
R639 vdd.t509 vdd.t507 84.656
R640 vdd.t510 vdd.t517 84.656
R641 vdd.t517 vdd.t512 84.656
R642 vdd.t512 vdd.t508 84.656
R643 vdd.t508 vdd.t515 84.656
R644 vdd.t515 vdd.t513 84.656
R645 vdd.t513 vdd.t518 84.656
R646 vdd.t518 vdd.t516 84.656
R647 vdd.t516 vdd.t511 84.656
R648 vdd.n390 vdd.t1 79.218
R649 vdd.n360 vdd.t110 77.822
R650 vdd.n383 vdd.n382 76.838
R651 vdd.n396 vdd.n395 76.775
R652 vdd.t255 vdd.t83 76.426
R653 vdd.n370 vdd.n369 74.564
R654 vdd.n342 vdd.t400 72.623
R655 vdd.n291 vdd.n290 72.477
R656 vdd.n395 vdd.t547 72.282
R657 vdd.t544 vdd.t531 70.381
R658 vdd.t556 vdd.t528 70.381
R659 vdd.t343 vdd.n373 69.089
R660 vdd.t557 vdd.n341 66.586
R661 vdd.n384 vdd.n383 61.94
R662 vdd.n385 vdd.n384 61.94
R663 vdd.n386 vdd.n385 61.94
R664 vdd.n387 vdd.n386 61.94
R665 vdd.n400 vdd.t551 61.066
R666 vdd.t453 vdd.t240 60.722
R667 vdd.n371 vdd.n370 59.964
R668 vdd.n372 vdd.n371 59.964
R669 vdd.n373 vdd.n372 59.964
R670 vdd.n389 vdd.t115 52.938
R671 vdd.n390 vdd.t264 51.299
R672 vdd.n585 vdd.t510 50.264
R673 vdd.n65 vdd.n59 49.509
R674 vdd.n598 vdd.t633 45.551
R675 vdd.n593 vdd.t642 45.551
R676 vdd.t547 vdd.t539 37.753
R677 vdd.n219 vdd.t142 37.605
R678 vdd.n341 vdd.t45 37.605
R679 vdd.n351 vdd.t392 37.26
R680 vdd.n363 vdd.n362 34.851
R681 vdd.n375 vdd.n363 34.851
R682 vdd.n228 vdd.t120 34.5
R683 vdd.t514 vdd.n585 34.391
R684 vdd.t264 vdd.t494 32.455
R685 vdd.n598 vdd.t606 29.329
R686 vdd.n599 vdd.t682 29.329
R687 vdd.n600 vdd.t628 29.329
R688 vdd.n601 vdd.t609 29.329
R689 vdd.n602 vdd.t648 29.329
R690 vdd.n597 vdd.t630 29.329
R691 vdd.n596 vdd.t601 29.329
R692 vdd.n595 vdd.t638 29.329
R693 vdd.n594 vdd.t623 29.329
R694 vdd.n593 vdd.t667 29.329
R695 vdd.t209 vdd.t64 28.29
R696 vdd.t64 vdd.t78 28.29
R697 vdd.t78 vdd.t172 28.29
R698 vdd.t172 vdd.t31 28.29
R699 vdd.t16 vdd.t11 28.29
R700 vdd.t250 vdd.t16 28.29
R701 vdd.t6 vdd.t250 28.29
R702 vdd.t331 vdd.t6 28.29
R703 vdd.t308 vdd.t331 28.29
R704 vdd.t291 vdd.t308 28.29
R705 vdd.t196 vdd.t291 28.29
R706 vdd.t177 vdd.t196 28.29
R707 vdd.t142 vdd.t177 28.29
R708 vdd.t120 vdd.t88 28.29
R709 vdd.t88 vdd.t55 28.29
R710 vdd.t55 vdd.t321 28.29
R711 vdd.t321 vdd.t40 28.29
R712 vdd.t40 vdd.t26 28.29
R713 vdd.t26 vdd.t286 28.29
R714 vdd.t245 vdd.t352 28.29
R715 vdd.t235 vdd.t245 28.29
R716 vdd.t326 vdd.t235 28.29
R717 vdd.t226 vdd.t326 28.29
R718 vdd.t281 vdd.t226 28.29
R719 vdd.t191 vdd.t281 28.29
R720 vdd.t525 vdd.t548 28.29
R721 vdd.t548 vdd.t519 28.29
R722 vdd.t519 vdd.t546 28.29
R723 vdd.t546 vdd.t543 28.29
R724 vdd.t543 vdd.t541 28.29
R725 vdd.t541 vdd.t535 28.29
R726 vdd.t506 vdd.t545 28.29
R727 vdd.t531 vdd.t506 28.29
R728 vdd.t550 vdd.t544 28.29
R729 vdd.t540 vdd.t550 28.29
R730 vdd.t536 vdd.t540 28.29
R731 vdd.t534 vdd.t536 28.29
R732 vdd.t526 vdd.t534 28.29
R733 vdd.t533 vdd.t532 28.29
R734 vdd.t532 vdd.t530 28.29
R735 vdd.t530 vdd.t556 28.29
R736 vdd.t528 vdd.t537 28.29
R737 vdd.t537 vdd.t505 28.29
R738 vdd.t524 vdd.t527 28.29
R739 vdd.t521 vdd.t524 28.29
R740 vdd.t554 vdd.t521 28.29
R741 vdd.t529 vdd.t554 28.29
R742 vdd.t553 vdd.t529 28.29
R743 vdd.t551 vdd.t553 28.29
R744 vdd.t523 vdd.t520 28.29
R745 vdd.t520 vdd.t522 28.29
R746 vdd.t522 vdd.t555 28.29
R747 vdd.t555 vdd.t552 28.29
R748 vdd.t552 vdd.t542 28.29
R749 vdd.t542 vdd.t549 28.29
R750 vdd.t114 vdd.t268 24.528
R751 vdd.t295 vdd.t114 24.528
R752 vdd.n290 vdd.t209 23.632
R753 vdd.n218 vdd.n217 23.406
R754 vdd.n399 vdd.t538 20.718
R755 vdd.n146 vdd.n145 19.059
R756 vdd.t268 vdd.n374 18.941
R757 vdd.n376 vdd.t276 18.933
R758 vdd.n102 vdd.n101 18.914
R759 vdd.n586 vdd.t514 18.518
R760 vdd.n71 vdd.n70 17.954
R761 vdd.n73 vdd.n72 17.254
R762 vdd.n74 vdd.n73 17.254
R763 vdd.n75 vdd.n74 17.254
R764 vdd.n76 vdd.n75 17.254
R765 vdd.n77 vdd.n76 17.254
R766 vdd.n78 vdd.n77 17.254
R767 vdd.n79 vdd.n78 17.254
R768 vdd.n68 vdd.n67 17.254
R769 vdd.n69 vdd.n68 17.254
R770 vdd.n70 vdd.n69 17.254
R771 vdd.n148 vdd.n147 17.254
R772 vdd.n149 vdd.n148 17.254
R773 vdd.n150 vdd.n149 17.254
R774 vdd.n139 vdd.n138 17.254
R775 vdd.n140 vdd.n139 17.254
R776 vdd.n141 vdd.n140 17.254
R777 vdd.n142 vdd.n141 17.254
R778 vdd.n143 vdd.n142 17.254
R779 vdd.n144 vdd.n143 17.254
R780 vdd.n145 vdd.n144 17.254
R781 vdd.n104 vdd.n103 17.254
R782 vdd.n105 vdd.n104 17.254
R783 vdd.n106 vdd.n105 17.254
R784 vdd.n95 vdd.n94 17.254
R785 vdd.n96 vdd.n95 17.254
R786 vdd.n97 vdd.n96 17.254
R787 vdd.n98 vdd.n97 17.254
R788 vdd.n99 vdd.n98 17.254
R789 vdd.n100 vdd.n99 17.254
R790 vdd.n101 vdd.n100 17.254
R791 vdd.n406 vdd.t397 17.25
R792 vdd.t115 vdd.t186 16.751
R793 vdd.n345 vdd.t375 16.387
R794 vdd.n594 vdd.n593 16.222
R795 vdd.n595 vdd.n594 16.222
R796 vdd.n596 vdd.n595 16.222
R797 vdd.n597 vdd.n596 16.222
R798 vdd.n602 vdd.n601 16.222
R799 vdd.n601 vdd.n600 16.222
R800 vdd.n600 vdd.n599 16.222
R801 vdd.n599 vdd.n598 16.222
R802 vdd.n403 vdd.t533 15.525
R803 vdd.n151 vdd.n150 14.308
R804 vdd.n107 vdd.n106 14.03
R805 vdd.t507 vdd.n589 13.756
R806 vdd.n410 vdd.t383 13.282
R807 vdd.n403 vdd.t526 12.765
R808 vdd.t549 vdd.n399 12.765
R809 vdd.n348 vdd.t407 12.42
R810 vdd.n362 vdd.t136 12.3
R811 vdd.t276 vdd.n375 12.3
R812 vdd.n362 vdd.t150 12.227
R813 vdd.n375 vdd.t295 12.227
R814 vdd.n80 vdd.n79 10.38
R815 vdd.n289 vdd.n288 10.062
R816 vdd.n400 vdd.t523 9.315
R817 vdd.t303 vdd.n376 9.168
R818 vdd.n374 vdd.t343 9.164
R819 vdd.n383 vdd.t263 9.125
R820 vdd.n384 vdd.t239 9.125
R821 vdd.n385 vdd.t167 9.125
R822 vdd.n386 vdd.t124 9.125
R823 vdd.n363 vdd.t82 9.125
R824 vdd.n363 vdd.t92 9.125
R825 vdd.n370 vdd.t299 9.125
R826 vdd.n371 vdd.t259 9.125
R827 vdd.n372 vdd.t217 9.125
R828 vdd.n373 vdd.t163 9.125
R829 vdd.n387 vdd.t303 9.125
R830 vdd.n319 vdd.n317 9.1
R831 vdd.n317 vdd.n135 9.1
R832 vdd.n262 vdd.n260 9.1
R833 vdd.n260 vdd.n258 9.1
R834 vdd.n258 vdd.n137 9.1
R835 vdd.t154 vdd.t312 8.174
R836 vdd.t200 vdd.t364 8.174
R837 vdd.n603 vdd.n597 8.111
R838 vdd.n603 vdd.n602 8.111
R839 vdd.n344 vdd.n1 7.03
R840 vdd vdd.n592 6.852
R841 vdd.t594 vdd.t137 6.63
R842 vdd.n398 vdd.n397 6.3
R843 vdd.n397 vdd.n396 6.3
R844 vdd.n408 vdd.n407 6.3
R845 vdd.n407 vdd.n406 6.3
R846 vdd.n402 vdd.n401 6.3
R847 vdd.n401 vdd.n400 6.3
R848 vdd.n347 vdd.n346 6.3
R849 vdd.n346 vdd.n345 6.3
R850 vdd.n350 vdd.n349 6.3
R851 vdd.n349 vdd.n348 6.3
R852 vdd.n357 vdd.n356 6.3
R853 vdd.n356 vdd.n355 6.3
R854 vdd.n412 vdd.n411 6.3
R855 vdd.n411 vdd.n410 6.3
R856 vdd.n344 vdd.n343 6.3
R857 vdd.n343 vdd.n342 6.3
R858 vdd.n492 vdd.n491 6.3
R859 vdd.n292 vdd.n289 5.95
R860 vdd.n49 vdd.n48 5.95
R861 vdd.n396 vdd.t155 5.932
R862 vdd.n288 vdd.n287 5.862
R863 vdd.n61 vdd.n60 5.862
R864 vdd.n461 vdd.n460 5.758
R865 vdd.n394 vdd.n393 5.192
R866 vdd.n353 vdd.n352 4.5
R867 vdd.n352 vdd.n351 4.5
R868 vdd.n415 vdd.n414 4.5
R869 vdd.n414 vdd.n413 4.5
R870 vdd.n409 vdd.n359 4.5
R871 vdd.n359 vdd.n358 4.5
R872 vdd.n490 vdd.n489 4.5
R873 vdd.n487 vdd.n486 4.355
R874 vdd.n388 vdd.n387 4.105
R875 vdd.n109 vdd.n107 4.004
R876 vdd.n232 vdd.n151 4
R877 vdd.n81 vdd.n80 4
R878 vdd vdd.n603 4
R879 vdd.n336 vdd.n57 3.725
R880 vdd.n335 vdd.n57 3.725
R881 vdd.n334 vdd.n56 3.725
R882 vdd.n333 vdd.n55 3.725
R883 vdd.n332 vdd.n54 3.725
R884 vdd.n331 vdd.n53 3.725
R885 vdd.n330 vdd.n51 3.725
R886 vdd.n215 vdd.n85 3.724
R887 vdd.n214 vdd.n86 3.724
R888 vdd.n213 vdd.n87 3.724
R889 vdd.n212 vdd.n88 3.724
R890 vdd.n211 vdd.n89 3.724
R891 vdd.n210 vdd.n90 3.724
R892 vdd.n209 vdd.n91 3.724
R893 vdd.n207 vdd.n93 3.724
R894 vdd.n340 vdd.n339 3.71
R895 vdd.n588 vdd.n587 3.626
R896 vdd.n338 vdd.n51 3.408
R897 vdd.n215 vdd.n84 3.4
R898 vdd.n207 vdd.n83 3.393
R899 vdd.n394 vdd.n361 3.15
R900 vdd.n361 vdd.n360 3.15
R901 vdd.n392 vdd.n391 3.15
R902 vdd.n391 vdd.n390 3.15
R903 vdd.n405 vdd.n404 3.15
R904 vdd.n404 vdd.n403 3.15
R905 vdd.n109 vdd.n108 3.15
R906 vdd.n112 vdd.n111 3.15
R907 vdd.n115 vdd.n114 3.15
R908 vdd.n114 vdd.n113 3.15
R909 vdd.n118 vdd.n117 3.15
R910 vdd.n117 vdd.n116 3.15
R911 vdd.n121 vdd.n120 3.15
R912 vdd.n120 vdd.n119 3.15
R913 vdd.n124 vdd.n123 3.15
R914 vdd.n123 vdd.n122 3.15
R915 vdd.n127 vdd.n126 3.15
R916 vdd.n126 vdd.n125 3.15
R917 vdd.n130 vdd.n129 3.15
R918 vdd.n129 vdd.n128 3.15
R919 vdd.n133 vdd.n132 3.15
R920 vdd.n132 vdd.n131 3.15
R921 vdd.n320 vdd.n319 3.15
R922 vdd.n319 vdd.n318 3.15
R923 vdd.n317 pmos_3p3_CDNS_679510442371_1.B 3.15
R924 vdd.n317 vdd.n316 3.15
R925 vdd.n315 vdd.n135 3.15
R926 vdd.n135 vdd.n134 3.15
R927 vdd.n314 vdd.n313 3.15
R928 vdd.n313 vdd.n312 3.15
R929 vdd.n311 vdd.n310 3.15
R930 vdd.n310 vdd.n309 3.15
R931 vdd.n308 vdd.n307 3.15
R932 vdd.n307 vdd.n306 3.15
R933 vdd.n305 vdd.n304 3.15
R934 vdd.n304 vdd.n303 3.15
R935 vdd.n302 vdd.n301 3.15
R936 vdd.n301 vdd.n300 3.15
R937 vdd.n299 vdd.n298 3.15
R938 vdd.n298 vdd.n297 3.15
R939 vdd.n296 vdd.n295 3.15
R940 vdd.n295 vdd.n294 3.15
R941 vdd.n293 vdd.n292 3.15
R942 vdd.n292 vdd.n291 3.15
R943 vdd.n287 vdd.n285 3.15
R944 vdd.n287 vdd.n286 3.15
R945 vdd.n284 vdd.n283 3.15
R946 vdd.n283 vdd.n282 3.15
R947 vdd.n281 vdd.n280 3.15
R948 vdd.n280 vdd.n279 3.15
R949 vdd.n278 vdd.n277 3.15
R950 vdd.n277 vdd.n276 3.15
R951 vdd.n275 vdd.n274 3.15
R952 vdd.n274 vdd.n273 3.15
R953 vdd.n272 vdd.n271 3.15
R954 vdd.n271 vdd.n270 3.15
R955 vdd.n269 vdd.n268 3.15
R956 vdd.n268 vdd.n267 3.15
R957 vdd.n266 vdd.n265 3.15
R958 vdd.n265 vdd.n264 3.15
R959 vdd.n263 vdd.n262 3.15
R960 vdd.n262 vdd.n261 3.15
R961 vdd.n260 pmos_3p3_CDNS_679510442370_1.B 3.15
R962 vdd.n260 vdd.n259 3.15
R963 vdd.n258 pmos_3p3_CDNS_679510442370_1.S 3.15
R964 vdd.n258 vdd.n257 3.15
R965 vdd.n256 vdd.n137 3.15
R966 vdd.n137 vdd.n136 3.15
R967 vdd.n255 vdd.n254 3.15
R968 vdd.n254 vdd.n253 3.15
R969 vdd.n252 vdd.n251 3.15
R970 vdd.n251 vdd.n250 3.15
R971 vdd.n249 vdd.n248 3.15
R972 vdd.n248 vdd.n247 3.15
R973 vdd.n246 vdd.n245 3.15
R974 vdd.n245 vdd.n244 3.15
R975 vdd.n243 vdd.n242 3.15
R976 vdd.n242 vdd.n241 3.15
R977 vdd.n240 vdd.n239 3.15
R978 vdd.n239 vdd.n238 3.15
R979 vdd.n237 vdd.n236 3.15
R980 vdd.n234 vdd.n233 3.15
R981 vdd.n203 vdd.n202 3.15
R982 vdd.n222 vdd.n221 3.15
R983 vdd.n154 vdd.n153 3.15
R984 vdd.n173 vdd.n172 3.15
R985 vdd.n176 vdd.n175 3.15
R986 vdd.n179 vdd.n178 3.15
R987 vdd.n182 vdd.n181 3.15
R988 vdd.n185 vdd.n184 3.15
R989 vdd.n188 vdd.n187 3.15
R990 vdd.n192 vdd.n191 3.15
R991 vdd.n224 vdd.n223 3.15
R992 vdd.n230 vdd.n229 3.15
R993 vdd.n229 vdd.n228 3.15
R994 vdd.n46 vdd.n45 3.15
R995 vdd.n41 vdd.n40 3.15
R996 vdd.n43 vdd.n42 3.15
R997 vdd.n36 vdd.n35 3.15
R998 vdd.n38 vdd.n37 3.15
R999 vdd.n31 vdd.n30 3.15
R1000 vdd.n33 vdd.n32 3.15
R1001 vdd.n24 vdd.n23 3.15
R1002 vdd.n28 vdd.n27 3.15
R1003 vdd.n26 vdd.n25 3.15
R1004 vdd.n21 vdd.n20 3.15
R1005 vdd.n16 vdd.n15 3.15
R1006 vdd.n18 vdd.n17 3.15
R1007 vdd.n11 vdd.n10 3.15
R1008 vdd.n13 vdd.n12 3.15
R1009 vdd.n6 vdd.n5 3.15
R1010 vdd.n8 vdd.n7 3.15
R1011 vdd.n3 vdd.n2 3.15
R1012 vdd.n226 vdd.n225 3.15
R1013 vdd.n62 vdd.n61 3.15
R1014 vdd.n204 vdd.n82 3.15
R1015 vdd.n219 vdd.n206 3.15
R1016 vdd.n341 vdd.n49 3.15
R1017 vdd.n341 vdd.n50 3.15
R1018 pmos_3p3_CDNS_679510442371_0.B vdd.n59 3.15
R1019 vdd.n66 vdd.n65 3.15
R1020 vdd.n65 vdd.n64 3.15
R1021 vdd.n219 vdd.n218 3.15
R1022 vdd.n219 vdd.n216 3.15
R1023 vdd.n589 vdd.n588 3.15
R1024 vdd.n587 vdd.n586 3.15
R1025 vdd.n585 vdd.n584 3.15
R1026 vdd.t509 vdd.n591 3.15
R1027 vdd.n408 vdd.n405 3.146
R1028 vdd.n230 vdd.n226 3.131
R1029 vdd.n64 vdd.t191 3.105
R1030 vdd.n170 vdd.n168 3.092
R1031 vdd.n377 vdd.t109 3.041
R1032 vdd.n378 vdd.t68 3.041
R1033 vdd.n379 vdd.t49 3.041
R1034 vdd.n380 vdd.t20 3.041
R1035 vdd.n381 vdd.t96 3.041
R1036 vdd.n382 vdd.t335 3.041
R1037 vdd.n364 vdd.t159 3.041
R1038 vdd.n365 vdd.t132 3.041
R1039 vdd.n366 vdd.t105 3.041
R1040 vdd.n367 vdd.t73 3.041
R1041 vdd.n368 vdd.t146 3.041
R1042 vdd.n369 vdd.t0 3.041
R1043 vdd.n582 vdd.n581 2.734
R1044 vdd.n405 vdd.n402 2.643
R1045 vdd.n162 vdd.n161 2.642
R1046 vdd.n191 vdd.n190 2.642
R1047 vdd.n187 vdd.n186 2.642
R1048 vdd.n184 vdd.n183 2.642
R1049 vdd.n181 vdd.n180 2.642
R1050 vdd.n178 vdd.n177 2.642
R1051 vdd.n175 vdd.n174 2.642
R1052 vdd.n172 vdd.n171 2.642
R1053 vdd.n153 vdd.n152 2.642
R1054 vdd.n166 vdd.n165 2.642
R1055 vdd.n164 vdd.n163 2.642
R1056 vdd.n162 vdd.n160 2.642
R1057 vdd.n158 vdd.n157 2.642
R1058 vdd.n156 vdd.n155 2.642
R1059 vdd.n190 vdd.n189 2.642
R1060 vdd.n449 vdd.n448 2.484
R1061 vdd.t494 vdd.t453 2.442
R1062 vdd.t561 vdd.t594 2.442
R1063 vdd.t186 vdd.t255 2.442
R1064 vdd.n80 vdd.n71 2.316
R1065 vdd.n592 vdd.n582 2.27
R1066 vdd.n592 vdd.t509 2.25
R1067 vdd.n503 vdd.n502 2.175
R1068 vdd.n402 vdd.n398 2.141
R1069 vdd.n327 pmos_3p3_CDNS_679510442370_0.D 2.062
R1070 vdd.n329 pmos_3p3_CDNS_679510442370_0.D 2.061
R1071 vdd.n324 pmos_3p3_CDNS_679510442370_0.D 2.061
R1072 vdd.n328 pmos_3p3_CDNS_679510442370_0.D 2.059
R1073 vdd.n326 pmos_3p3_CDNS_679510442370_0.D 2.059
R1074 vdd.n325 pmos_3p3_CDNS_679510442370_0.D 2.059
R1075 vdd.n323 pmos_3p3_CDNS_679510442370_0.D 2.059
R1076 vdd.n322 pmos_3p3_CDNS_679510442370_0.D 2.057
R1077 vdd.t509 vdd.n590 2.011
R1078 vdd.n44 vdd.n41 1.863
R1079 vdd.n39 vdd.n36 1.863
R1080 vdd.n34 vdd.n31 1.863
R1081 vdd.n29 vdd.n24 1.863
R1082 vdd.n25 vdd.n22 1.863
R1083 vdd.n19 vdd.n16 1.863
R1084 vdd.n14 vdd.n11 1.863
R1085 vdd.n9 vdd.n6 1.863
R1086 vdd.n4 vdd.n3 1.863
R1087 vdd.n225 vdd.n4 1.862
R1088 vdd.n9 vdd.n8 1.862
R1089 vdd.n14 vdd.n13 1.862
R1090 vdd.n19 vdd.n18 1.862
R1091 vdd.n22 vdd.n21 1.862
R1092 vdd.n29 vdd.n28 1.862
R1093 vdd.n34 vdd.n33 1.862
R1094 vdd.n39 vdd.n38 1.862
R1095 vdd.n44 vdd.n43 1.862
R1096 vdd.n47 vdd.n46 1.855
R1097 vdd.n61 vdd.n47 1.855
R1098 vdd.n340 vdd.n59 1.855
R1099 vdd.n219 vdd.n156 1.83
R1100 vdd.n219 vdd.n158 1.83
R1101 vdd.n219 vdd.n159 1.83
R1102 vdd.n219 vdd.n162 1.83
R1103 vdd.n219 vdd.n164 1.83
R1104 vdd.n219 vdd.n166 1.83
R1105 vdd.n219 vdd.n167 1.83
R1106 vdd.n376 vdd.t254 1.75
R1107 vdd.n546 vdd.n545 1.704
R1108 vdd.n554 vdd 1.558
R1109 vdd.n170 vdd.n169 1.546
R1110 vdd.n337 vdd.n49 1.546
R1111 vdd.n221 vdd.n220 1.546
R1112 vdd.n374 vdd.t185 1.544
R1113 vdd.n534 vdd.n533 1.538
R1114 vdd.n218 vdd.n92 1.533
R1115 vdd.n205 vdd.n203 1.519
R1116 vdd.n205 vdd.n204 1.519
R1117 vdd.n501 vdd.n500 1.503
R1118 vdd.n525 vdd.n524 1.503
R1119 vdd.n416 vdd.n415 1.501
R1120 vdd.n354 vdd.n353 1.5
R1121 vdd.n151 vdd.n146 1.488
R1122 vdd.n531 vdd.n495 1.461
R1123 vdd.n107 vdd.n102 1.365
R1124 vdd.n480 vdd.n479 1.333
R1125 vdd.n229 vdd.n227 1.288
R1126 vdd.n518 vdd.n517 1.26
R1127 vdd.n543 vdd.n542 1.126
R1128 vdd.n494 vdd.n493 1.125
R1129 vdd.n581 vdd.n421 1.124
R1130 vdd.n438 vdd.n437 1.121
R1131 vdd.n547 vdd.n546 1.121
R1132 vdd.n580 vdd.n579 1.121
R1133 vdd.n445 vdd.n444 1.121
R1134 vdd.n464 vdd.n463 1.121
R1135 vdd.n472 vdd.n471 1.121
R1136 vdd.n458 vdd.n457 1.121
R1137 vdd.n474 vdd.n473 1.121
R1138 vdd.n447 vdd.n446 1.12
R1139 vdd.n460 vdd.n459 1.12
R1140 vdd.n524 vdd.n523 1.102
R1141 vdd.n536 vdd.n481 1.092
R1142 vdd.n508 vdd.n507 1.084
R1143 pmos_3p3_CDNS_679510442371_0.B vdd.n92 1.079
R1144 pmos_3p3_CDNS_679510442371_0.B vdd.n84 1.075
R1145 vdd.n219 vdd.n170 1.071
R1146 vdd.n220 vdd.n219 1.07
R1147 pmos_3p3_CDNS_679510442371_0.B vdd.n337 1.07
R1148 pmos_3p3_CDNS_679510442371_0.B vdd.n338 1.07
R1149 vdd.n393 vdd.n389 0.939
R1150 vdd.n515 vdd.n514 0.861
R1151 vdd.n219 vdd.n205 0.817
R1152 pmos_3p3_CDNS_679510442371_0.B vdd.n83 0.811
R1153 vdd.n543 vdd.n475 0.718
R1154 vdd.n539 vdd.n538 0.696
R1155 vdd.n493 vdd.n485 0.677
R1156 vdd.n529 vdd.n528 0.65
R1157 vdd.n341 vdd.n47 0.649
R1158 vdd.n339 pmos_3p3_CDNS_679510442371_0.B 0.649
R1159 vdd.n341 vdd.n340 0.649
R1160 vdd.n341 vdd.n44 0.645
R1161 vdd.n341 vdd.n39 0.645
R1162 vdd.n341 vdd.n34 0.645
R1163 vdd.n341 vdd.n29 0.645
R1164 vdd.n341 vdd.n22 0.645
R1165 vdd.n341 vdd.n19 0.645
R1166 vdd.n341 vdd.n14 0.645
R1167 vdd.n341 vdd.n9 0.645
R1168 vdd.n341 vdd.n4 0.645
R1169 vdd.n341 vdd.n58 0.645
R1170 pmos_3p3_CDNS_679510442371_0.B vdd.n336 0.645
R1171 vdd.n341 vdd.n57 0.645
R1172 pmos_3p3_CDNS_679510442371_0.B vdd.n335 0.645
R1173 vdd.n341 vdd.n56 0.645
R1174 pmos_3p3_CDNS_679510442371_0.B vdd.n334 0.645
R1175 vdd.n341 vdd.n55 0.645
R1176 pmos_3p3_CDNS_679510442371_0.B vdd.n333 0.645
R1177 vdd.n341 vdd.n54 0.645
R1178 pmos_3p3_CDNS_679510442371_0.B vdd.n332 0.645
R1179 vdd.n341 vdd.n53 0.645
R1180 pmos_3p3_CDNS_679510442371_0.B vdd.n331 0.645
R1181 vdd.n341 vdd.n52 0.645
R1182 pmos_3p3_CDNS_679510442371_0.B vdd.n330 0.645
R1183 vdd.n341 vdd.n51 0.645
R1184 pmos_3p3_CDNS_679510442371_0.B vdd.n91 0.645
R1185 pmos_3p3_CDNS_679510442371_0.B vdd.n90 0.645
R1186 pmos_3p3_CDNS_679510442371_0.B vdd.n89 0.645
R1187 pmos_3p3_CDNS_679510442371_0.B vdd.n88 0.645
R1188 pmos_3p3_CDNS_679510442371_0.B vdd.n87 0.645
R1189 pmos_3p3_CDNS_679510442371_0.B vdd.n86 0.645
R1190 pmos_3p3_CDNS_679510442371_0.B vdd.n85 0.645
R1191 pmos_3p3_CDNS_679510442371_0.B vdd.n93 0.645
R1192 vdd.n219 vdd.n208 0.645
R1193 vdd.n219 vdd.n209 0.645
R1194 vdd.n219 vdd.n210 0.645
R1195 vdd.n219 vdd.n211 0.645
R1196 vdd.n219 vdd.n212 0.645
R1197 vdd.n219 vdd.n213 0.645
R1198 vdd.n219 vdd.n214 0.645
R1199 vdd.n219 vdd.n215 0.645
R1200 vdd.n219 vdd.n207 0.645
R1201 vdd.n511 vdd.n510 0.634
R1202 vdd.n398 vdd.n394 0.502
R1203 vdd.n409 vdd.n408 0.399
R1204 vdd.n231 vdd.n224 0.356
R1205 vdd.n329 vdd.n63 0.325
R1206 vdd.n582 vdd.n0 0.318
R1207 vdd.n329 vdd.n328 0.315
R1208 vdd.n328 vdd.n327 0.315
R1209 vdd.n327 vdd.n326 0.315
R1210 vdd.n325 vdd.n324 0.315
R1211 vdd.n324 vdd.n323 0.315
R1212 vdd.n323 vdd.n322 0.315
R1213 vdd vdd.n553 0.286
R1214 pmos_3p3_CDNS_679510442370_0.B vdd.n325 0.257
R1215 vdd.n111 vdd.n110 0.245
R1216 vdd.n236 vdd.n235 0.245
R1217 vdd.n418 vdd.n417 0.226
R1218 pmos_3p3_CDNS_679510442371_0.D vdd.n329 0.178
R1219 vdd.n328 pmos_3p3_CDNS_679510442371_0.D 0.178
R1220 vdd.n327 pmos_3p3_CDNS_679510442371_0.D 0.178
R1221 vdd.n326 pmos_3p3_CDNS_679510442371_0.D 0.178
R1222 vdd.n325 pmos_3p3_CDNS_679510442371_0.D 0.178
R1223 vdd.n324 pmos_3p3_CDNS_679510442371_0.D 0.178
R1224 vdd.n323 pmos_3p3_CDNS_679510442371_0.D 0.178
R1225 vdd.n322 pmos_3p3_CDNS_679510442371_0.D 0.178
R1226 vdd.n500 vdd.n499 0.176
R1227 vdd.n481 vdd.n478 0.152
R1228 pmos_3p3_CDNS_679510442371_0.B vdd.n63 0.143
R1229 pmos_3p3_CDNS_679510442370_1.B vdd.n82 0.141
R1230 vdd.n495 vdd.n484 0.136
R1231 vdd.n201 vdd.n200 0.13
R1232 vdd.n200 vdd.n199 0.13
R1233 vdd.n199 vdd.n198 0.13
R1234 vdd.n198 vdd.n197 0.13
R1235 vdd.n197 vdd.n196 0.13
R1236 vdd.n196 vdd.n195 0.13
R1237 vdd.n195 vdd.n194 0.13
R1238 vdd.n194 vdd.n193 0.13
R1239 vdd.n192 vdd.n188 0.13
R1240 vdd.n188 vdd.n185 0.13
R1241 vdd.n185 vdd.n182 0.13
R1242 vdd.n182 vdd.n179 0.13
R1243 vdd.n179 vdd.n176 0.13
R1244 vdd.n176 vdd.n173 0.13
R1245 vdd.n173 vdd.n154 0.13
R1246 vdd.n222 vdd.n154 0.13
R1247 vdd.n224 vdd.n222 0.13
R1248 vdd.n202 vdd.n201 0.128
R1249 pmos_3p3_CDNS_679510442370_0.B vdd.n192 0.128
R1250 pmos_3p3_CDNS_679510442370_0.B vdd.n26 0.128
R1251 vdd.n322 vdd.n82 0.125
R1252 vdd.n232 vdd.n231 0.121
R1253 vdd.n514 vdd.n512 0.116
R1254 vdd.n493 vdd.n492 0.105
R1255 vdd.n524 vdd.n522 0.104
R1256 vdd.n522 vdd.n521 0.102
R1257 vdd.n507 vdd.n505 0.099
R1258 vdd.n492 vdd.n490 0.098
R1259 vdd.n393 vdd.n392 0.094
R1260 vdd.n507 vdd.n506 0.086
R1261 vdd.n63 vdd.n62 0.083
R1262 vdd.n353 vdd.n350 0.082
R1263 vdd.n495 vdd.n494 0.069
R1264 vdd.n514 vdd.n513 0.068
R1265 vdd.n350 vdd.n347 0.06
R1266 vdd.n326 pmos_3p3_CDNS_679510442370_0.B 0.057
R1267 vdd.n481 vdd.n480 0.052
R1268 vdd.n389 vdd.n388 0.047
R1269 vdd.n542 vdd.n541 0.042
R1270 vdd.n483 vdd.n482 0.022
R1271 vdd.n541 vdd.n540 0.021
R1272 vdd.n231 vdd.n230 0.018
R1273 vdd.n488 vdd.n487 0.018
R1274 vdd.n551 vdd.n550 0.017
R1275 vdd.n432 vdd.n431 0.016
R1276 vdd.n437 vdd.n435 0.016
R1277 vdd.n428 vdd.n427 0.015
R1278 vdd.n347 vdd.n344 0.015
R1279 vdd.n415 vdd.n357 0.015
R1280 vdd.n415 vdd.n412 0.015
R1281 vdd.n412 vdd.n409 0.015
R1282 vdd.n499 vdd.n498 0.014
R1283 vdd.n545 vdd.n544 0.014
R1284 vdd.n450 vdd.n449 0.014
R1285 vdd.n437 vdd.n436 0.014
R1286 vdd.n455 vdd.n454 0.013
R1287 vdd.n447 vdd.n434 0.013
R1288 vdd.n558 vdd.n557 0.012
R1289 vdd.n471 vdd.n470 0.012
R1290 vdd.n448 vdd.n447 0.012
R1291 vdd.n463 vdd.n462 0.012
R1292 vdd.n427 vdd.n426 0.012
R1293 vdd.n426 vdd.n425 0.012
R1294 vdd.n459 vdd.n433 0.012
R1295 vdd.n459 vdd.n458 0.012
R1296 vdd.n552 vdd.n551 0.012
R1297 vdd.n477 vdd.n476 0.011
R1298 vdd.n474 vdd.n429 0.011
R1299 vdd.n475 vdd.n474 0.011
R1300 vdd.n540 vdd.n539 0.011
R1301 vdd.n425 vdd.n424 0.01
R1302 vdd.n424 vdd.n423 0.01
R1303 vdd.n453 vdd.n452 0.01
R1304 vdd.n457 vdd.n453 0.01
R1305 vdd.n473 vdd.n464 0.01
R1306 vdd.n473 vdd.n472 0.01
R1307 vdd.n468 vdd.n467 0.01
R1308 vdd.n467 vdd.n466 0.01
R1309 vdd.n464 vdd.n461 0.01
R1310 vdd.n469 vdd.n468 0.01
R1311 vdd.n472 vdd.n469 0.01
R1312 vdd.n466 vdd.n465 0.01
R1313 vdd.n457 vdd.n456 0.01
R1314 vdd.n452 vdd.n451 0.01
R1315 vdd.n446 vdd.n438 0.01
R1316 vdd.n438 vdd.n0 0.009
R1317 vdd.n441 vdd.n440 0.009
R1318 vdd.n442 vdd.n441 0.009
R1319 vdd.n445 vdd.n443 0.009
R1320 vdd.n581 vdd.n580 0.009
R1321 vdd.n576 vdd.n575 0.009
R1322 vdd.n574 vdd.n573 0.009
R1323 vdd.n572 vdd.n571 0.009
R1324 vdd.n570 vdd.n569 0.009
R1325 vdd.n568 vdd.n567 0.009
R1326 vdd.n566 vdd.n565 0.009
R1327 vdd.n564 vdd.n563 0.009
R1328 vdd.n562 vdd.n561 0.009
R1329 vdd.n560 vdd.n559 0.009
R1330 vdd.n556 vdd.n555 0.009
R1331 vdd.n549 vdd.n548 0.009
R1332 vdd.n548 vdd.n547 0.009
R1333 vdd.n443 vdd.n442 0.009
R1334 vdd.n547 vdd.n422 0.009
R1335 vdd.n555 vdd.n554 0.009
R1336 vdd.n559 vdd.n558 0.009
R1337 vdd.n563 vdd.n562 0.009
R1338 vdd.n567 vdd.n566 0.009
R1339 vdd.n571 vdd.n570 0.009
R1340 vdd.n575 vdd.n574 0.009
R1341 vdd.n550 vdd.n549 0.009
R1342 vdd.n573 vdd.n572 0.009
R1343 vdd.n569 vdd.n568 0.009
R1344 vdd.n565 vdd.n564 0.009
R1345 vdd.n561 vdd.n560 0.009
R1346 vdd.n580 vdd.n576 0.009
R1347 vdd.n440 vdd.n439 0.009
R1348 vdd.n446 vdd.n445 0.009
R1349 vdd.n433 vdd.n432 0.008
R1350 vdd.n546 vdd.n428 0.008
R1351 vdd.n520 vdd.n519 0.008
R1352 vdd.n544 vdd.n543 0.007
R1353 vdd.n458 vdd.n450 0.007
R1354 vdd.n456 vdd.n455 0.007
R1355 vdd.n460 vdd.n430 0.007
R1356 vdd.n557 vdd.n556 0.006
R1357 vdd.n553 vdd.n552 0.006
R1358 pmos_3p3_CDNS_679510442370_1.B pmos_3p3_CDNS_679510442371_1.B 0.006
R1359 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1360 pmos_3p3_CDNS_679510442371_0.S pmos_3p3_CDNS_679510442371_0.D 0.005
R1361 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1362 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1363 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1364 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1365 pmos_3p3_CDNS_679510442371_0.S pmos_3p3_CDNS_679510442371_0.D 0.005
R1366 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1367 pmos_3p3_CDNS_679510442371_0.S pmos_3p3_CDNS_679510442371_0.D 0.005
R1368 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.S 0.005
R1369 pmos_3p3_CDNS_679510442371_0.S pmos_3p3_CDNS_679510442371_0.D 0.005
R1370 vdd.n421 vdd.n418 0.004
R1371 vdd.n234 vdd.n232 0.004
R1372 pmos_3p3_CDNS_679510442371_0.B vdd.n321 0.004
R1373 pmos_3p3_CDNS_679510442371_0.D pmos_3p3_CDNS_679510442371_0.B 0.004
R1374 pmos_3p3_CDNS_679510442371_0.D vdd.n1 0.004
R1375 pmos_3p3_CDNS_679510442371_0.S vdd.n81 0.004
R1376 pmos_3p3_CDNS_679510442371_0.B pmos_3p3_CDNS_679510442371_0.S 0.004
R1377 vdd.n515 vdd.n511 0.004
R1378 vdd.n421 vdd.n420 0.004
R1379 vdd.n535 vdd.n534 0.003
R1380 vdd.n525 vdd.n518 0.003
R1381 vdd.n502 vdd.n501 0.003
R1382 vdd.n112 vdd.n109 0.003
R1383 vdd.n115 vdd.n112 0.003
R1384 vdd.n118 vdd.n115 0.003
R1385 vdd.n121 vdd.n118 0.003
R1386 vdd.n124 vdd.n121 0.003
R1387 vdd.n127 vdd.n124 0.003
R1388 vdd.n130 vdd.n127 0.003
R1389 vdd.n133 vdd.n130 0.003
R1390 pmos_3p3_CDNS_679510442371_1.B vdd.n315 0.003
R1391 vdd.n315 vdd.n314 0.003
R1392 vdd.n314 vdd.n311 0.003
R1393 vdd.n311 vdd.n308 0.003
R1394 vdd.n308 vdd.n305 0.003
R1395 vdd.n305 vdd.n302 0.003
R1396 vdd.n302 vdd.n299 0.003
R1397 vdd.n299 vdd.n296 0.003
R1398 vdd.n296 vdd.n293 0.003
R1399 vdd.n293 pmos_3p3_CDNS_679510442371_1.B 0.003
R1400 vdd.n285 pmos_3p3_CDNS_679510442370_1.B 0.003
R1401 vdd.n285 vdd.n284 0.003
R1402 vdd.n284 vdd.n281 0.003
R1403 vdd.n281 vdd.n278 0.003
R1404 vdd.n278 vdd.n275 0.003
R1405 vdd.n275 vdd.n272 0.003
R1406 vdd.n272 vdd.n269 0.003
R1407 vdd.n269 vdd.n266 0.003
R1408 vdd.n266 vdd.n263 0.003
R1409 vdd.n263 pmos_3p3_CDNS_679510442370_1.B 0.003
R1410 pmos_3p3_CDNS_679510442370_1.S vdd.n256 0.003
R1411 vdd.n256 vdd.n255 0.003
R1412 vdd.n255 vdd.n252 0.003
R1413 vdd.n252 vdd.n249 0.003
R1414 vdd.n249 vdd.n246 0.003
R1415 vdd.n246 vdd.n243 0.003
R1416 vdd.n243 vdd.n240 0.003
R1417 vdd.n240 vdd.n237 0.003
R1418 vdd.n237 vdd.n234 0.003
R1419 pmos_3p3_CDNS_679510442371_0.S vdd.n66 0.003
R1420 vdd.n579 vdd.n578 0.003
R1421 vdd.n578 vdd.n577 0.003
R1422 vdd.n508 vdd.n504 0.002
R1423 vdd.n510 vdd.n509 0.002
R1424 vdd.n517 vdd.n516 0.002
R1425 vdd.n538 vdd.n537 0.002
R1426 vdd.n537 vdd.n536 0.002
R1427 vdd.n516 vdd.n515 0.002
R1428 vdd.n504 vdd.n503 0.002
R1429 vdd.n509 vdd.n508 0.002
R1430 vdd.n420 vdd.n419 0.002
R1431 vdd.n532 vdd.n531 0.002
R1432 pmos_3p3_CDNS_679510442371_1.B pmos_3p3_CDNS_679510442371_1.S 0.002
R1433 pmos_3p3_CDNS_679510442370_1.S pmos_3p3_CDNS_679510442370_1.B 0.002
R1434 pmos_3p3_CDNS_679510442371_0.S pmos_3p3_CDNS_679510442371_0.B 0.002
R1435 pmos_3p3_CDNS_679510442371_0.B pmos_3p3_CDNS_679510442371_0.D 0.002
R1436 pmos_3p3_CDNS_679510442371_0.D vdd.n66 0.002
R1437 vdd.n533 vdd.n532 0.002
R1438 vdd.n501 vdd.n497 0.002
R1439 vdd.n526 vdd.n525 0.002
R1440 vdd.n536 vdd.n535 0.002
R1441 vdd.n497 vdd.n496 0.002
R1442 vdd.n321 vdd.n133 0.001
R1443 vdd.n321 vdd.n320 0.001
R1444 vdd.n320 pmos_3p3_CDNS_679510442371_1.S 0.001
R1445 vdd.n193 pmos_3p3_CDNS_679510442370_0.B 0.001
R1446 vdd.n27 pmos_3p3_CDNS_679510442370_0.B 0.001
R1447 pmos_3p3_CDNS_679510442371_0.S vdd.n1 0.001
R1448 vdd.n81 pmos_3p3_CDNS_679510442371_0.D 0.001
R1449 vdd.n521 vdd.n520 0.001
R1450 vdd.n490 vdd.n488 0.001
R1451 vdd.n484 vdd.n483 0.001
R1452 vdd.n478 vdd.n477 0.001
R1453 vdd.n416 vdd.n354 0.001
R1454 vdd.n417 vdd.n416 0.001
R1455 vdd.n528 vdd.n527 0.001
R1456 vdd.n530 vdd.n529 0.001
R1457 vdd.n531 vdd.n530 0.001
R1458 vdd.n527 vdd.n526 0.001
R1459 vin1.n83 vin1.n82 298.834
R1460 vin1.n74 vin1.t15 166.643
R1461 vin1.n65 vin1.t61 166.643
R1462 vin1.n76 vin1.t9 156.018
R1463 vin1.n68 vin1.t25 153.907
R1464 vin1.n69 vin1.t28 153.907
R1465 vin1.n71 vin1.t20 153.907
R1466 vin1.n80 vin1.t69 153.907
R1467 vin1.n74 vin1.t30 153.907
R1468 vin1.n75 vin1.t32 153.907
R1469 vin1.n77 vin1.t26 153.907
R1470 vin1.n78 vin1.t2 153.907
R1471 vin1.n79 vin1.t77 153.907
R1472 vin1.n81 vin1.t71 153.907
R1473 vin1.n82 vin1.t64 153.907
R1474 vin1.n73 vin1.t49 153.907
R1475 vin1.n72 vin1.t44 153.907
R1476 vin1.n70 vin1.t36 153.907
R1477 vin1.n67 vin1.t17 153.907
R1478 vin1.n66 vin1.t76 153.907
R1479 vin1.n65 vin1.t11 153.907
R1480 vin1.n35 vin1.t57 151.863
R1481 vin1.n10 vin1.t70 151.854
R1482 vin1.n46 vin1.t12 149.61
R1483 vin1.n0 vin1.t56 147.42
R1484 vin1.n64 vin1.t27 136.874
R1485 vin1.n63 vin1.t13 136.874
R1486 vin1.n62 vin1.t37 136.874
R1487 vin1.n61 vin1.t40 136.874
R1488 vin1.n60 vin1.t45 136.874
R1489 vin1.n59 vin1.t68 136.874
R1490 vin1.n58 vin1.t48 136.874
R1491 vin1.n57 vin1.t51 136.874
R1492 vin1.n56 vin1.t53 136.874
R1493 vin1.n55 vin1.t4 136.874
R1494 vin1.n54 vin1.t58 136.874
R1495 vin1.n53 vin1.t39 136.874
R1496 vin1.n52 vin1.t43 136.874
R1497 vin1.n51 vin1.t66 136.874
R1498 vin1.n50 vin1.t75 136.874
R1499 vin1.n49 vin1.t0 136.874
R1500 vin1.n48 vin1.t5 136.874
R1501 vin1.n47 vin1.t55 136.874
R1502 vin1.n46 vin1.t7 136.874
R1503 vin1.n35 vin1.t41 135.901
R1504 vin1.n36 vin1.t74 135.901
R1505 vin1.n37 vin1.t47 135.901
R1506 vin1.n38 vin1.t34 135.901
R1507 vin1.n39 vin1.t8 135.901
R1508 vin1.n40 vin1.t62 135.901
R1509 vin1.n41 vin1.t18 135.901
R1510 vin1.n42 vin1.t72 135.901
R1511 vin1.n43 vin1.t50 135.901
R1512 vin1.n18 vin1.t1 135.901
R1513 vin1.n17 vin1.t31 135.901
R1514 vin1.n16 vin1.t6 135.901
R1515 vin1.n15 vin1.t73 135.901
R1516 vin1.n14 vin1.t46 135.901
R1517 vin1.n13 vin1.t79 135.901
R1518 vin1.n12 vin1.t54 135.901
R1519 vin1.n11 vin1.t29 135.901
R1520 vin1.n10 vin1.t60 135.901
R1521 vin1.n34 vin1.t10 135.901
R1522 vin1.n33 vin1.t65 135.901
R1523 vin1.n32 vin1.t42 135.901
R1524 vin1.n31 vin1.t21 135.901
R1525 vin1.n30 vin1.t59 135.901
R1526 vin1.n29 vin1.t35 135.901
R1527 vin1.n28 vin1.t14 135.901
R1528 vin1.n27 vin1.t63 135.901
R1529 vin1.n26 vin1.t19 135.901
R1530 vin1.n25 vin1.t3 135.901
R1531 vin1.n8 vin1.t24 134.684
R1532 vin1.n7 vin1.t78 134.684
R1533 vin1.n6 vin1.t38 134.684
R1534 vin1.n5 vin1.t16 134.684
R1535 vin1.n4 vin1.t67 134.684
R1536 vin1.n3 vin1.t23 134.684
R1537 vin1.n2 vin1.t22 134.684
R1538 vin1.n1 vin1.t52 134.684
R1539 vin1.n0 vin1.t33 134.684
R1540 vin1.n44 vin1.n34 44.082
R1541 vin1.n44 vin1.n43 43.179
R1542 vin1.n25 vin1.n24 43.176
R1543 vin1.n19 vin1.n18 32.801
R1544 vin1.n55 vin1.n54 31.685
R1545 vin1.n9 vin1.n8 25.765
R1546 vin1.n83 vin1.n73 25.472
R1547 vin1.n36 vin1.n35 15.962
R1548 vin1.n37 vin1.n36 15.962
R1549 vin1.n38 vin1.n37 15.962
R1550 vin1.n39 vin1.n38 15.962
R1551 vin1.n40 vin1.n39 15.962
R1552 vin1.n41 vin1.n40 15.962
R1553 vin1.n42 vin1.n41 15.962
R1554 vin1.n43 vin1.n42 15.962
R1555 vin1.n18 vin1.n17 15.962
R1556 vin1.n17 vin1.n16 15.962
R1557 vin1.n16 vin1.n15 15.962
R1558 vin1.n15 vin1.n14 15.962
R1559 vin1.n14 vin1.n13 15.962
R1560 vin1.n13 vin1.n12 15.962
R1561 vin1.n12 vin1.n11 15.962
R1562 vin1.n11 vin1.n10 15.962
R1563 vin1.n34 vin1.n33 15.962
R1564 vin1.n33 vin1.n32 15.962
R1565 vin1.n32 vin1.n31 15.962
R1566 vin1.n31 vin1.n30 15.962
R1567 vin1.n30 vin1.n29 15.962
R1568 vin1.n29 vin1.n28 15.962
R1569 vin1.n28 vin1.n27 15.962
R1570 vin1.n27 vin1.n26 15.962
R1571 vin1.n26 vin1.n25 15.962
R1572 vin1 vin1.n87 15.635
R1573 vin1.n85 vin1.n84 13.151
R1574 vin1.n77 vin1.n76 12.891
R1575 vin1.n8 vin1.n7 12.736
R1576 vin1.n7 vin1.n6 12.736
R1577 vin1.n6 vin1.n5 12.736
R1578 vin1.n5 vin1.n4 12.736
R1579 vin1.n4 vin1.n3 12.736
R1580 vin1.n3 vin1.n2 12.736
R1581 vin1.n2 vin1.n1 12.736
R1582 vin1.n1 vin1.n0 12.736
R1583 vin1.n64 vin1.n63 12.736
R1584 vin1.n63 vin1.n62 12.736
R1585 vin1.n62 vin1.n61 12.736
R1586 vin1.n61 vin1.n60 12.736
R1587 vin1.n60 vin1.n59 12.736
R1588 vin1.n59 vin1.n58 12.736
R1589 vin1.n58 vin1.n57 12.736
R1590 vin1.n57 vin1.n56 12.736
R1591 vin1.n56 vin1.n55 12.736
R1592 vin1.n54 vin1.n53 12.736
R1593 vin1.n53 vin1.n52 12.736
R1594 vin1.n52 vin1.n51 12.736
R1595 vin1.n51 vin1.n50 12.736
R1596 vin1.n50 vin1.n49 12.736
R1597 vin1.n49 vin1.n48 12.736
R1598 vin1.n48 vin1.n47 12.736
R1599 vin1.n47 vin1.n46 12.736
R1600 vin1.n66 vin1.n65 12.736
R1601 vin1.n67 vin1.n66 12.736
R1602 vin1.n68 vin1.n67 12.736
R1603 vin1.n69 vin1.n68 12.736
R1604 vin1.n70 vin1.n69 12.736
R1605 vin1.n71 vin1.n70 12.736
R1606 vin1.n72 vin1.n71 12.736
R1607 vin1.n73 vin1.n72 12.736
R1608 vin1.n82 vin1.n81 12.736
R1609 vin1.n81 vin1.n80 12.736
R1610 vin1.n80 vin1.n79 12.736
R1611 vin1.n79 vin1.n78 12.736
R1612 vin1.n78 vin1.n77 12.736
R1613 vin1.n75 vin1.n74 12.736
R1614 vin1.n76 vin1.n75 12.58
R1615 vin1.n86 vin1.n44 12.065
R1616 vin1.n84 vin1.n83 10.39
R1617 vin1.n84 vin1.n64 9.834
R1618 vin1.n21 vin1.n20 1.5
R1619 vin1.n86 vin1.n85 1.498
R1620 vin1.n24 vin1.n23 1.123
R1621 vin1.n20 vin1.n19 0.039
R1622 vin1.n86 vin1.n9 0.03
R1623 vin1.n87 vin1.n86 0.017
R1624 vin1.n85 vin1.n45 0.01
R1625 vin1.n23 vin1.n22 0.009
R1626 vin1.n22 vin1.n21 0.005
R1627 vout_t.n15 vout_t.n0 35.786
R1628 vout_t.n0 vout_t 6.794
R1629 vout_t.n12 vout_t.n1 4.5
R1630 vout_t.n11 vout_t.n10 4.5
R1631 vout_t.n16 vout_t.n15 3.135
R1632 vout_t.n15 vout_t.n14 2.38
R1633 vout_t.n13 vout_t.n7 2.358
R1634 vout_t.n8 vout_t.n7 2.253
R1635 vout_t.n14 vout_t.n13 0.897
R1636 vout_t.n9 vout_t.n8 0.897
R1637 vout_t.n5 vout_t.n4 0.626
R1638 vout_t.n4 nmos_3p3_CDNS_679510442372_0.D 0.626
R1639 nmos_3p3_CDNS_679510442372_0.D vout_t.n3 0.626
R1640 vout_t.n3 vout_t.n2 0.626
R1641 vout_t.n18 vout_t.n17 0.626
R1642 vout_t vout_t.n18 0.626
R1643 vout_t vout_t.n20 0.626
R1644 vout_t.n20 vout_t.n19 0.626
R1645 vout_t.n9 vout_t.n0 0.592
R1646 vout_t.n16 vout_t 0.478
R1647 vout_t.n17 vout_t 0.477
R1648 vout_t.n18 vout_t 0.477
R1649 vout_t.n20 vout_t 0.477
R1650 vout_t.n19 vout_t 0.477
R1651 vout_t.n6 nmos_3p3_CDNS_679510442372_0.D 0.313
R1652 nmos_3p3_CDNS_679510442372_0.D vout_t.n5 0.313
R1653 vout_t.n2 nmos_3p3_CDNS_679510442372_0.D 0.313
R1654 vout_t vout_t.n16 0.313
R1655 vout_t.n17 vout_t 0.313
R1656 vout_t.n19 vout_t 0.313
R1657 vout_t.n7 vout_t.n6 0.299
R1658 vout_t.n6 nmos_3p3_CDNS_679510442372_0.D 0.285
R1659 vout_t.n5 nmos_3p3_CDNS_679510442372_0.D 0.285
R1660 vout_t.n4 nmos_3p3_CDNS_679510442372_0.D 0.285
R1661 vout_t.n3 nmos_3p3_CDNS_679510442372_0.D 0.285
R1662 vout_t.n2 nmos_3p3_CDNS_679510442372_0.D 0.285
R1663 vout_t.n10 vout_t.n1 0.068
R1664 vout_t.n12 vout_t.n11 0.063
R1665 vout_t.n10 vout_t.n9 0.032
R1666 vout_t.n14 vout_t.n1 0.032
R1667 vout_t.n13 vout_t.n12 0.024
R1668 vout_t.n11 vout_t.n8 0.024
R1669 vbiasp vbiasp.t5 69.282
R1670 vbiasp.n3 vbiasp.n2 36.278
R1671 vbiasp.n2 vbiasp.n1 24.078
R1672 vbiasp.n3 vbiasp.n0 24.078
R1673 vbiasp.n3 vbiasp.t6 12.166
R1674 vbiasp.n1 vbiasp.t4 12.166
R1675 vbiasp.n1 vbiasp.t2 12.166
R1676 vbiasp.n2 vbiasp.t0 12.166
R1677 vbiasp.n2 vbiasp.t7 12.166
R1678 vbiasp.n0 vbiasp.t3 12.166
R1679 vbiasp.n0 vbiasp.t1 12.166
R1680 vbiasp.t5 vbiasp.n3 12.166
R1681 vprog vprog.t0 16.77
R1682 vbiasn.n2 vbiasn.t0 58.837
R1683 vbiasn.n0 vbiasn.t3 58.837
R1684 vbiasn.n4 vbiasn.n2 46.64
R1685 vbiasn.n2 vbiasn.t2 36.5
R1686 vbiasn.n0 vbiasn.t1 36.5
R1687 vbiasn.n1 vbiasn.n0 33.863
R1688 vbiasn vbiasn.n8 28.211
R1689 vbiasn.n5 vbiasn.n4 2.244
R1690 vbiasn.n5 vbiasn.n1 0.756
R1691 vbiasn.n7 vbiasn.n6 0.024
R1692 vbiasn.n4 vbiasn.n3 0.015
R1693 vbiasn.n8 vbiasn.n7 0.005
R1694 vbiasn.n6 vbiasn.n5 0.002
C0 vin1 vbiasp 0.19fF
C1 vin2 vdd 12.39fF
C2 a_9856_n4071# vin1 8.71fF
C3 vin1 a_4788_4131# 0.04fF
C4 a_19749_n6676# a_7580_3503# 0.36fF
C5 a_35590_n7073# vbiasn 0.00fF
C6 vbiasn a_19749_n2296# 0.01fF
C7 vbiasp vbiasn 4.77fF
C8 vin1 a_21261_4878# 0.00fF
C9 vbiasn a_4788_4131# 3.46fF
C10 vin1 a_7580_3503# 3.97fF
C11 vdd a_13786_2835# 2.35fF
C12 vbiasn a_21261_4878# 0.08fF
C13 vdd a_13786_5007# 7.45fF
C14 vdd a_6084_4175# 3.51fF
C15 vbiasn a_5010_6963# 0.05fF
C16 vout a_13786_2835# 5.40fF
C17 vdd a_5796_4175# 0.48fF
C18 vout a_13786_5007# 2.00fF
C19 a_9656_n5262# a_5884_4131# 0.01fF
C20 vdd a_4700_4175# 2.87fF
C21 vin2 a_13786_2835# 7.96fF
C22 a_11072_n909# a_5884_4131# 0.05fF
C23 vin2 a_13786_5007# 1.00fF
C24 vprog vdd 3.09fF
C25 a_28902_5067# vout_t 0.01fF
C26 vin2 a_6084_4175# 1.43fF
C27 a_35590_n7073# vdd 0.23fF
C28 a_19749_n2296# vdd 8.97fF
C29 vbiasp vdd 7.63fF
C30 a_9856_n4071# vdd 4.31fF
C31 a_4788_4131# vdd 3.87fF
C32 a_13786_5007# a_13786_2835# 3.94fF
C33 a_11072_n909# a_9656_n5262# 0.08fF
C34 a_11312_n4152# a_9656_n5262# 0.33fF
C35 a_11512_n3371# vdd 0.22fF
C36 a_21261_4878# vdd 26.48fF
C37 a_35590_n7073# vout 0.23fF
C38 a_11312_n4152# a_11072_n909# 0.01fF
C39 a_19749_n2296# vout 0.00fF
C40 vbiasp vout 0.01fF
C41 a_7580_3503# vdd 17.47fF
C42 a_4788_4131# vout 0.01fF
C43 a_5010_6963# vdd 2.83fF
C44 vin2 a_19749_n2296# 0.43fF
C45 vin2 vbiasp 0.31fF
C46 a_21261_4878# vout 1.51fF
C47 a_9856_n4071# vin2 6.59fF
C48 a_5796_5519# vdd 40.42fF
C49 vin2 a_4788_4131# 4.07fF
C50 a_5796_4175# a_6084_4175# 0.81fF
C51 a_31806_5067# a_31806_2835# 2.36fF
C52 vbiasn a_5884_4131# 0.09fF
C53 vin2 a_21261_4878# 0.20fF
C54 a_4700_4175# a_6084_4175# 0.00fF
C55 a_28902_5067# a_31806_2835# 3.87fF
C56 a_19749_n2296# a_13786_2835# 0.07fF
C57 vbiasp a_13786_2835# 5.64fF
C58 vin1 a_9656_n5262# 0.06fF
C59 vin2 a_7580_3503# 4.17fF
C60 a_4700_4175# a_5796_4175# 0.01fF
C61 a_28902_5067# a_31806_5067# 0.37fF
C62 a_19749_n6676# a_31806_2835# 0.00fF
C63 a_4788_4131# a_13786_2835# 0.07fF
C64 a_19749_n2296# a_13786_5007# 0.46fF
C65 vbiasp a_13786_5007# 0.50fF
C66 vin2 a_5010_6963# 0.12fF
C67 a_19749_n6676# a_31806_5067# 0.02fF
C68 a_35590_n7073# a_6084_4175# 0.00fF
C69 a_4788_4131# a_13786_5007# 0.04fF
C70 a_21261_4878# a_13786_2835# 0.03fF
C71 vbiasp a_6084_4175# 1.41fF
C72 vin2 a_5796_5519# 0.00fF
C73 a_19749_n6676# a_28902_5067# 2.09fF
C74 a_9856_n4071# a_6084_4175# 0.04fF
C75 a_7580_3503# a_13786_2835# 30.08fF
C76 a_21261_4878# a_13786_5007# 0.54fF
C77 a_4788_4131# a_6084_4175# 0.19fF
C78 a_11512_n3371# a_6084_4175# 0.60fF
C79 a_31806_2835# vbiasn 1.24fF
C80 a_7580_3503# a_13786_5007# 30.08fF
C81 a_4788_4131# a_5796_4175# 0.19fF
C82 a_21261_4878# a_6084_4175# 0.50fF
C83 vbiasp a_4700_4175# 0.01fF
C84 vdd vout_t 2.10fF
C85 a_31806_5067# vbiasn 1.53fF
C86 a_7580_3503# a_6084_4175# 0.02fF
C87 a_4788_4131# a_4700_4175# 1.01fF
C88 vin1 a_19749_n6676# 0.72fF
C89 a_28902_5067# vbiasn 0.29fF
C90 a_5010_6963# a_6084_4175# 0.19fF
C91 a_5796_5519# a_13786_5007# 0.00fF
C92 vprog a_4788_4131# 0.00fF
C93 vbiasp a_19749_n2296# 2.86fF
C94 a_19749_n6676# vbiasn 0.06fF
C95 a_5796_5519# a_6084_4175# 0.36fF
C96 vdd a_5884_4131# 4.55fF
C97 vout_t vout 4.31fF
C98 a_9856_n4071# a_19749_n2296# 27.21fF
C99 a_4788_4131# a_19749_n2296# 0.08fF
C100 vbiasp a_4788_4131# 0.08fF
C101 a_5010_6963# a_4700_4175# 0.33fF
C102 a_5796_5519# a_5796_4175# 0.60fF
C103 a_35590_n7073# a_21261_4878# 0.25fF
C104 a_9856_n4071# a_4788_4131# 0.98fF
C105 a_21261_4878# a_19749_n2296# 6.97fF
C106 vin1 vbiasn 0.04fF
C107 vbiasp a_21261_4878# 2.82fF
C108 a_11512_n3371# a_9856_n4071# 0.18fF
C109 a_5796_5519# a_4700_4175# 0.01fF
C110 vprog a_5010_6963# 0.12fF
C111 a_11512_n3371# a_4788_4131# 0.71fF
C112 a_7580_3503# a_19749_n2296# 0.42fF
C113 a_21261_4878# a_4788_4131# 0.28fF
C114 vbiasp a_7580_3503# 0.15fF
C115 a_9656_n5262# vdd 0.40fF
C116 vprog a_5796_5519# 0.11fF
C117 a_7580_3503# a_4788_4131# 0.00fF
C118 vbiasp a_5010_6963# 0.06fF
C119 a_11072_n909# vdd 0.17fF
C120 vin2 a_5884_4131# 0.10fF
C121 a_9856_n4071# a_5010_6963# 0.80fF
C122 a_11312_n4152# vdd 0.28fF
C123 a_7580_3503# a_21261_4878# 0.00fF
C124 a_5010_6963# a_4788_4131# 2.30fF
C125 vbiasp a_5796_5519# 0.01fF
C126 a_31806_2835# vdd 1.42fF
C127 a_11512_n3371# a_5010_6963# 0.53fF
C128 a_5796_5519# a_4788_4131# 0.60fF
C129 a_31806_5067# vdd 6.33fF
C130 a_28902_5067# vdd 7.66fF
C131 a_5796_5519# a_7580_3503# 4.49fF
C132 a_31806_2835# vout 24.04fF
C133 a_19749_n6676# vdd 5.92fF
C134 a_5796_5519# a_5010_6963# 0.06fF
C135 a_31806_5067# vout 0.43fF
C136 a_5884_4131# a_6084_4175# 0.80fF
C137 a_28902_5067# vout 19.95fF
C138 a_5884_4131# a_5796_4175# 0.33fF
C139 vin1 vdd 17.25fF
C140 a_19749_n6676# vout 0.00fF
C141 vbiasn vdd 1.42fF
C142 a_31806_2835# a_13786_2835# 0.89fF
C143 a_19749_n6676# vin2 3.56fF
C144 a_11072_n909# a_6084_4175# 0.11fF
C145 a_31806_5067# a_13786_2835# 0.44fF
C146 a_31806_2835# a_13786_5007# 0.04fF
C147 a_11312_n4152# a_6084_4175# 0.90fF
C148 vbiasp a_5884_4131# 0.09fF
C149 a_31806_5067# a_13786_5007# 0.97fF
C150 a_28902_5067# a_13786_2835# 0.20fF
C151 a_31806_2835# a_6084_4175# 0.45fF
C152 vin1 vin2 3.60fF
C153 a_9856_n4071# a_5884_4131# 0.00fF
C154 vbiasn vout 0.14fF
C155 a_4788_4131# a_5884_4131# 0.08fF
C156 a_28902_5067# a_13786_5007# 0.23fF
C157 a_31806_5067# a_6084_4175# 0.33fF
C158 a_19749_n6676# a_13786_2835# 0.03fF
C159 vin2 vbiasn 0.56fF
C160 a_19749_n6676# a_13786_5007# 0.05fF
C161 a_28902_5067# a_6084_4175# 0.58fF
C162 a_7580_3503# a_5884_4131# 0.21fF
C163 vin1 a_13786_2835# 1.54fF
C164 a_19749_n6676# a_6084_4175# 0.01fF
C165 a_9856_n4071# a_9656_n5262# 3.76fF
C166 a_5010_6963# a_5884_4131# 0.07fF
C167 a_9656_n5262# a_4788_4131# 0.00fF
C168 vin1 a_13786_5007# 6.54fF
C169 a_11512_n3371# a_9656_n5262# 0.25fF
C170 a_9856_n4071# a_11072_n909# 0.07fF
C171 a_35590_n7073# a_31806_2835# 0.02fF
C172 a_11312_n4152# a_9856_n4071# 0.22fF
C173 vbiasn a_13786_2835# 1.32fF
C174 a_5796_5519# a_5884_4131# 2.87fF
C175 a_11072_n909# a_4788_4131# 0.01fF
C176 vin1 a_6084_4175# 0.07fF
C177 a_31806_2835# vbiasp 0.00fF
C178 a_11312_n4152# a_4788_4131# 0.42fF
C179 a_11512_n3371# a_11072_n909# 0.07fF
C180 vbiasn a_13786_5007# 0.45fF
C181 a_11312_n4152# a_11512_n3371# 0.53fF
C182 a_31806_5067# a_19749_n2296# 0.01fF
C183 a_31806_2835# a_4788_4131# 0.36fF
C184 a_31806_5067# vbiasp 0.04fF
C185 vbiasn a_6084_4175# 0.15fF
C186 a_31806_5067# a_4788_4131# 0.30fF
C187 a_28902_5067# a_19749_n2296# 1.44fF
C188 a_9656_n5262# a_5010_6963# 3.12fF
C189 a_31806_2835# a_21261_4878# 0.05fF
C190 a_28902_5067# vbiasp 2.11fF
C191 a_28902_5067# a_4788_4131# 0.39fF
C192 a_31806_5067# a_21261_4878# 0.59fF
C193 a_19749_n6676# a_19749_n2296# 6.61fF
C194 a_11072_n909# a_5010_6963# 0.06fF
C195 a_19749_n6676# vbiasp 2.40fF
C196 a_11312_n4152# a_5010_6963# 0.02fF
C197 a_9856_n4071# a_19749_n6676# 27.39fF
C198 vdd vout 13.56fF
C199 a_28902_5067# a_21261_4878# 1.74fF
C200 a_19749_n6676# a_4788_4131# 0.09fF
C201 vin1 a_19749_n2296# 3.55fF
C202 a_19749_n6676# a_21261_4878# 5.31fF
C203 vbiasn vss 7.78fF
C204 vbiasp vss 9.49fF
C205 vin2 vss 25.62fF
C206 vin1 vss 31.23fF
C207 vprog vss 2.10fF
C208 a_35590_n7073# vss 2.29fF $ **FLOATING
C209 a_9856_n4071# vss 4.41fF
C210 a_11512_n3371# vss 0.23fF
C211 a_11312_n4152# vss 1.33fF
C212 a_9656_n5262# vss 15.02fF
C213 a_11072_n909# vss 1.01fF
C214 a_31806_2835# vss 25.35fF
C215 a_31806_5067# vss -3.14fF
C216 a_28902_5067# vss 22.67fF
C217 a_19749_n6676# vss 4.83fF
C218 a_13786_2835# vss -3.56fF
C219 a_13786_5007# vss -4.95fF
C220 a_6084_4175# vss 12.91fF
C221 a_5796_4175# vss -0.29fF
C222 a_4700_4175# vss -1.18fF
C223 a_5884_4131# vss -0.29fF
C224 a_19749_n2296# vss 2.03fF
C225 a_4788_4131# vss 1.34fF
C226 a_21261_4878# vss -2.74fF
C227 a_7580_3503# vss -4.63fF
C228 a_5010_6963# vss 6.31fF
C229 a_5796_5519# vss -2.21fF
C230 vout vss 21.72fF
C231 vout_t vss 6.82fF
C232 vdd vss 743.01fF
C233 vbiasn.t1 vss 0.27fF
C234 vbiasn.t3 vss 0.32fF
C235 vbiasn.n0 vss 0.20fF $ **FLOATING
C236 vbiasn.n1 vss 0.04fF $ **FLOATING
C237 vbiasn.t2 vss 0.27fF
C238 vbiasn.t0 vss 0.32fF
C239 vbiasn.n2 vss 0.21fF $ **FLOATING
C240 vbiasn.n3 vss 0.01fF $ **FLOATING
C241 vbiasn.n4 vss 0.18fF $ **FLOATING
C242 vbiasn.n5 vss 0.00fF $ **FLOATING
C243 vbiasn.n6 vss 0.00fF $ **FLOATING
C244 vbiasn.n7 vss 0.00fF $ **FLOATING
C245 vbiasn.n8 vss 3.52fF $ **FLOATING
C246 vprog.t0 vss 1.69fF
C247 vbiasp.t6 vss 1.47fF
C248 vbiasp.t3 vss 1.47fF
C249 vbiasp.t1 vss 1.47fF
C250 vbiasp.n0 vss 1.25fF $ **FLOATING
C251 vbiasp.t0 vss 1.47fF
C252 vbiasp.t7 vss 1.47fF
C253 vbiasp.t4 vss 1.47fF
C254 vbiasp.t2 vss 1.47fF
C255 vbiasp.n1 vss 1.25fF $ **FLOATING
C256 vbiasp.n2 vss 1.30fF $ **FLOATING
C257 vbiasp.n3 vss 1.30fF $ **FLOATING
C258 vbiasp.t5 vss 2.73fF
C259 vout_t.n0 vss 2.33fF $ **FLOATING
C260 vout_t.n1 vss 0.02fF $ **FLOATING
C261 nmos_3p3_CDNS_679510442372_0.D vss 0.70fF $ **FLOATING
C262 vout_t.n2 vss 0.06fF $ **FLOATING
C263 vout_t.n3 vss 0.07fF $ **FLOATING
C264 vout_t.n4 vss 0.07fF $ **FLOATING
C265 vout_t.n5 vss 0.06fF $ **FLOATING
C266 vout_t.n6 vss 0.05fF $ **FLOATING
C267 vout_t.n7 vss 0.07fF $ **FLOATING
C268 vout_t.n8 vss 0.02fF $ **FLOATING
C269 vout_t.n9 vss 0.10fF $ **FLOATING
C270 vout_t.n10 vss 0.02fF $ **FLOATING
C271 vout_t.n11 vss 0.02fF $ **FLOATING
C272 vout_t.n12 vss 0.02fF $ **FLOATING
C273 vout_t.n13 vss 0.02fF $ **FLOATING
C274 vout_t.n14 vss 0.37fF $ **FLOATING
C275 vout_t.n15 vss 1.07fF $ **FLOATING
C276 vout_t.n16 vss 0.42fF $ **FLOATING
C277 vout_t.n17 vss 0.08fF $ **FLOATING
C278 vout_t.n18 vss 0.10fF $ **FLOATING
C279 vout_t.n19 vss 0.08fF $ **FLOATING
C280 vout_t.n20 vss 0.10fF $ **FLOATING
C281 vin1.t24 vss 0.28fF
C282 vin1.t78 vss 0.28fF
C283 vin1.t38 vss 0.28fF
C284 vin1.t16 vss 0.28fF
C285 vin1.t67 vss 0.28fF
C286 vin1.t23 vss 0.28fF
C287 vin1.t22 vss 0.28fF
C288 vin1.t52 vss 0.28fF
C289 vin1.t33 vss 0.28fF
C290 vin1.t56 vss 0.29fF
C291 vin1.n0 vss 0.27fF $ **FLOATING
C292 vin1.n1 vss 0.15fF $ **FLOATING
C293 vin1.n2 vss 0.15fF $ **FLOATING
C294 vin1.n3 vss 0.15fF $ **FLOATING
C295 vin1.n4 vss 0.15fF $ **FLOATING
C296 vin1.n5 vss 0.15fF $ **FLOATING
C297 vin1.n6 vss 0.15fF $ **FLOATING
C298 vin1.n7 vss 0.15fF $ **FLOATING
C299 vin1.n8 vss 0.18fF $ **FLOATING
C300 vin1.n9 vss 0.27fF $ **FLOATING
C301 vin1.t10 vss 0.28fF
C302 vin1.t65 vss 0.28fF
C303 vin1.t42 vss 0.28fF
C304 vin1.t21 vss 0.28fF
C305 vin1.t59 vss 0.28fF
C306 vin1.t35 vss 0.28fF
C307 vin1.t14 vss 0.28fF
C308 vin1.t63 vss 0.28fF
C309 vin1.t19 vss 0.28fF
C310 vin1.t3 vss 0.28fF
C311 vin1.t1 vss 0.28fF
C312 vin1.t31 vss 0.28fF
C313 vin1.t6 vss 0.28fF
C314 vin1.t73 vss 0.28fF
C315 vin1.t46 vss 0.28fF
C316 vin1.t79 vss 0.28fF
C317 vin1.t54 vss 0.28fF
C318 vin1.t29 vss 0.28fF
C319 vin1.t60 vss 0.28fF
C320 vin1.t70 vss 0.29fF
C321 vin1.n10 vss 0.26fF $ **FLOATING
C322 vin1.n11 vss 0.14fF $ **FLOATING
C323 vin1.n12 vss 0.14fF $ **FLOATING
C324 vin1.n13 vss 0.14fF $ **FLOATING
C325 vin1.n14 vss 0.14fF $ **FLOATING
C326 vin1.n15 vss 0.14fF $ **FLOATING
C327 vin1.n16 vss 0.14fF $ **FLOATING
C328 vin1.n17 vss 0.14fF $ **FLOATING
C329 vin1.n18 vss 0.19fF $ **FLOATING
C330 vin1.n19 vss 0.46fF $ **FLOATING
C331 vin1.n20 vss 0.01fF $ **FLOATING
C332 vin1.n21 vss 0.01fF $ **FLOATING
C333 vin1.n22 vss 0.01fF $ **FLOATING
C334 vin1.n23 vss 0.01fF $ **FLOATING
C335 vin1.n24 vss 0.14fF $ **FLOATING
C336 vin1.n25 vss 0.17fF $ **FLOATING
C337 vin1.n26 vss 0.14fF $ **FLOATING
C338 vin1.n27 vss 0.14fF $ **FLOATING
C339 vin1.n28 vss 0.14fF $ **FLOATING
C340 vin1.n29 vss 0.14fF $ **FLOATING
C341 vin1.n30 vss 0.14fF $ **FLOATING
C342 vin1.n31 vss 0.14fF $ **FLOATING
C343 vin1.n32 vss 0.14fF $ **FLOATING
C344 vin1.n33 vss 0.14fF $ **FLOATING
C345 vin1.n34 vss 0.40fF $ **FLOATING
C346 vin1.t50 vss 0.28fF
C347 vin1.t72 vss 0.28fF
C348 vin1.t18 vss 0.28fF
C349 vin1.t62 vss 0.28fF
C350 vin1.t8 vss 0.28fF
C351 vin1.t34 vss 0.28fF
C352 vin1.t47 vss 0.28fF
C353 vin1.t74 vss 0.28fF
C354 vin1.t41 vss 0.28fF
C355 vin1.t57 vss 0.29fF
C356 vin1.n35 vss 0.26fF $ **FLOATING
C357 vin1.n36 vss 0.14fF $ **FLOATING
C358 vin1.n37 vss 0.14fF $ **FLOATING
C359 vin1.n38 vss 0.14fF $ **FLOATING
C360 vin1.n39 vss 0.14fF $ **FLOATING
C361 vin1.n40 vss 0.14fF $ **FLOATING
C362 vin1.n41 vss 0.14fF $ **FLOATING
C363 vin1.n42 vss 0.14fF $ **FLOATING
C364 vin1.n43 vss 0.17fF $ **FLOATING
C365 vin1.n44 vss 4.14fF $ **FLOATING
C366 vin1.n45 vss 0.06fF $ **FLOATING
C367 vin1.t27 vss 0.28fF
C368 vin1.t13 vss 0.28fF
C369 vin1.t37 vss 0.28fF
C370 vin1.t40 vss 0.28fF
C371 vin1.t45 vss 0.28fF
C372 vin1.t68 vss 0.28fF
C373 vin1.t48 vss 0.28fF
C374 vin1.t51 vss 0.28fF
C375 vin1.t53 vss 0.28fF
C376 vin1.t4 vss 0.28fF
C377 vin1.t58 vss 0.28fF
C378 vin1.t39 vss 0.28fF
C379 vin1.t43 vss 0.28fF
C380 vin1.t66 vss 0.28fF
C381 vin1.t75 vss 0.28fF
C382 vin1.t0 vss 0.28fF
C383 vin1.t5 vss 0.28fF
C384 vin1.t55 vss 0.28fF
C385 vin1.t7 vss 0.28fF
C386 vin1.t12 vss 0.29fF
C387 vin1.n46 vss 0.28fF $ **FLOATING
C388 vin1.n47 vss 0.15fF $ **FLOATING
C389 vin1.n48 vss 0.15fF $ **FLOATING
C390 vin1.n49 vss 0.15fF $ **FLOATING
C391 vin1.n50 vss 0.15fF $ **FLOATING
C392 vin1.n51 vss 0.15fF $ **FLOATING
C393 vin1.n52 vss 0.15fF $ **FLOATING
C394 vin1.n53 vss 0.15fF $ **FLOATING
C395 vin1.n54 vss 0.19fF $ **FLOATING
C396 vin1.n55 vss 0.19fF $ **FLOATING
C397 vin1.n56 vss 0.15fF $ **FLOATING
C398 vin1.n57 vss 0.15fF $ **FLOATING
C399 vin1.n58 vss 0.15fF $ **FLOATING
C400 vin1.n59 vss 0.15fF $ **FLOATING
C401 vin1.n60 vss 0.15fF $ **FLOATING
C402 vin1.n61 vss 0.15fF $ **FLOATING
C403 vin1.n62 vss 0.15fF $ **FLOATING
C404 vin1.n63 vss 0.15fF $ **FLOATING
C405 vin1.n64 vss 0.15fF $ **FLOATING
C406 vin1.t49 vss 0.29fF
C407 vin1.t44 vss 0.29fF
C408 vin1.t20 vss 0.29fF
C409 vin1.t36 vss 0.29fF
C410 vin1.t28 vss 0.29fF
C411 vin1.t25 vss 0.29fF
C412 vin1.t17 vss 0.29fF
C413 vin1.t76 vss 0.29fF
C414 vin1.t11 vss 0.29fF
C415 vin1.t61 vss 0.30fF
C416 vin1.n65 vss 0.30fF $ **FLOATING
C417 vin1.n66 vss 0.16fF $ **FLOATING
C418 vin1.n67 vss 0.16fF $ **FLOATING
C419 vin1.n68 vss 0.16fF $ **FLOATING
C420 vin1.n69 vss 0.16fF $ **FLOATING
C421 vin1.n70 vss 0.16fF $ **FLOATING
C422 vin1.n71 vss 0.16fF $ **FLOATING
C423 vin1.n72 vss 0.16fF $ **FLOATING
C424 vin1.n73 vss 0.19fF $ **FLOATING
C425 vin1.t64 vss 0.29fF
C426 vin1.t71 vss 0.29fF
C427 vin1.t69 vss 0.29fF
C428 vin1.t77 vss 0.29fF
C429 vin1.t2 vss 0.29fF
C430 vin1.t26 vss 0.29fF
C431 vin1.t9 vss 0.29fF
C432 vin1.t32 vss 0.29fF
C433 vin1.t30 vss 0.29fF
C434 vin1.t15 vss 0.30fF
C435 vin1.n74 vss 0.30fF $ **FLOATING
C436 vin1.n75 vss 0.16fF $ **FLOATING
C437 vin1.n76 vss 0.16fF $ **FLOATING
C438 vin1.n77 vss 0.16fF $ **FLOATING
C439 vin1.n78 vss 0.16fF $ **FLOATING
C440 vin1.n79 vss 0.16fF $ **FLOATING
C441 vin1.n80 vss 0.16fF $ **FLOATING
C442 vin1.n81 vss 0.16fF $ **FLOATING
C443 vin1.n82 vss 0.70fF $ **FLOATING
C444 vin1.n83 vss 0.94fF $ **FLOATING
C445 vin1.n84 vss 1.49fF $ **FLOATING
C446 vin1.n85 vss 0.98fF $ **FLOATING
C447 vin1.n86 vss 2.68fF $ **FLOATING
C448 vin1.n87 vss 5.64fF $ **FLOATING
C449 vdd.t509 vss 13.44fF
C450 vdd.n0 vss 3.34fF $ **FLOATING
C451 vdd.n1 vss 1.37fF $ **FLOATING
C452 vdd.t45 vss 1.62fF
C453 vdd.n2 vss 0.01fF $ **FLOATING
C454 vdd.n3 vss 0.01fF $ **FLOATING
C455 vdd.n5 vss 0.01fF $ **FLOATING
C456 vdd.n6 vss 0.01fF $ **FLOATING
C457 vdd.n7 vss 0.01fF $ **FLOATING
C458 vdd.n8 vss 0.01fF $ **FLOATING
C459 vdd.n10 vss 0.01fF $ **FLOATING
C460 vdd.n11 vss 0.01fF $ **FLOATING
C461 vdd.n12 vss 0.01fF $ **FLOATING
C462 vdd.n13 vss 0.01fF $ **FLOATING
C463 vdd.n15 vss 0.01fF $ **FLOATING
C464 vdd.n16 vss 0.01fF $ **FLOATING
C465 vdd.n17 vss 0.01fF $ **FLOATING
C466 vdd.n18 vss 0.01fF $ **FLOATING
C467 vdd.n20 vss 0.01fF $ **FLOATING
C468 vdd.n21 vss 0.01fF $ **FLOATING
C469 vdd.n23 vss 0.01fF $ **FLOATING
C470 vdd.n24 vss 0.01fF $ **FLOATING
C471 vdd.n25 vss 0.01fF $ **FLOATING
C472 vdd.n26 vss 0.01fF $ **FLOATING
C473 pmos_3p3_CDNS_679510442370_0.B vss 0.03fF $ **FLOATING
C474 vdd.n27 vss 0.01fF $ **FLOATING
C475 vdd.n28 vss 0.01fF $ **FLOATING
C476 vdd.n30 vss 0.01fF $ **FLOATING
C477 vdd.n31 vss 0.01fF $ **FLOATING
C478 vdd.n32 vss 0.01fF $ **FLOATING
C479 vdd.n33 vss 0.01fF $ **FLOATING
C480 vdd.n35 vss 0.01fF $ **FLOATING
C481 vdd.n36 vss 0.01fF $ **FLOATING
C482 vdd.n37 vss 0.01fF $ **FLOATING
C483 vdd.n38 vss 0.01fF $ **FLOATING
C484 vdd.n40 vss 0.01fF $ **FLOATING
C485 vdd.n41 vss 0.01fF $ **FLOATING
C486 vdd.n42 vss 0.01fF $ **FLOATING
C487 vdd.n43 vss 0.01fF $ **FLOATING
C488 vdd.n45 vss 0.01fF $ **FLOATING
C489 vdd.n46 vss 0.01fF $ **FLOATING
C490 vdd.n48 vss 0.17fF $ **FLOATING
C491 vdd.n49 vss 0.01fF $ **FLOATING
C492 vdd.n50 vss 0.01fF $ **FLOATING
C493 vdd.n51 vss 0.01fF $ **FLOATING
C494 vdd.n52 vss 0.01fF $ **FLOATING
C495 vdd.n53 vss 0.01fF $ **FLOATING
C496 vdd.n54 vss 0.01fF $ **FLOATING
C497 vdd.n55 vss 0.01fF $ **FLOATING
C498 vdd.n56 vss 0.01fF $ **FLOATING
C499 vdd.n57 vss 0.01fF $ **FLOATING
C500 vdd.n58 vss 0.01fF $ **FLOATING
C501 vdd.n59 vss 0.04fF $ **FLOATING
C502 vdd.n60 vss 0.16fF $ **FLOATING
C503 vdd.n61 vss 0.01fF $ **FLOATING
C504 vdd.n62 vss 0.01fF $ **FLOATING
C505 vdd.n63 vss 0.03fF $ **FLOATING
C506 vdd.t352 vss 1.46fF
C507 vdd.t245 vss 1.46fF
C508 vdd.t235 vss 1.46fF
C509 vdd.t326 vss 1.46fF
C510 vdd.t226 vss 1.46fF
C511 vdd.t281 vss 1.46fF
C512 vdd.t191 vss 0.81fF
C513 vdd.n64 vss 0.73fF $ **FLOATING
C514 vdd.n65 vss 0.21fF $ **FLOATING
C515 vdd.n66 vss 0.31fF $ **FLOATING
C516 pmos_3p3_CDNS_679510442370_0.D vss 3.37fF $ **FLOATING
C517 pmos_3p3_CDNS_679510442371_0.S vss 6.81fF $ **FLOATING
C518 pmos_3p3_CDNS_679510442371_0.D vss 6.87fF $ **FLOATING
C519 pmos_3p3_CDNS_679510442371_0.B vss 1.18fF $ **FLOATING
C520 vdd.t119 vss 0.14fF
C521 vdd.t87 vss 0.14fF
C522 vdd.n67 vss 0.11fF $ **FLOATING
C523 vdd.t54 vss 0.14fF
C524 vdd.n68 vss 0.06fF $ **FLOATING
C525 vdd.t320 vss 0.14fF
C526 vdd.n69 vss 0.06fF $ **FLOATING
C527 vdd.t39 vss 0.14fF
C528 vdd.n70 vss 0.06fF $ **FLOATING
C529 vdd.t25 vss 0.14fF
C530 vdd.n71 vss 0.06fF $ **FLOATING
C531 vdd.t44 vss 0.14fF
C532 vdd.t190 vss 0.14fF
C533 vdd.n72 vss 0.11fF $ **FLOATING
C534 vdd.t280 vss 0.14fF
C535 vdd.n73 vss 0.06fF $ **FLOATING
C536 vdd.t225 vss 0.14fF
C537 vdd.n74 vss 0.06fF $ **FLOATING
C538 vdd.t325 vss 0.14fF
C539 vdd.n75 vss 0.06fF $ **FLOATING
C540 vdd.t234 vss 0.14fF
C541 vdd.n76 vss 0.06fF $ **FLOATING
C542 vdd.t244 vss 0.14fF
C543 vdd.n77 vss 0.06fF $ **FLOATING
C544 vdd.t351 vss 0.14fF
C545 vdd.n78 vss 0.06fF $ **FLOATING
C546 vdd.t285 vss 0.14fF
C547 vdd.n79 vss 0.06fF $ **FLOATING
C548 vdd.n80 vss 0.01fF $ **FLOATING
C549 vdd.n81 vss 0.31fF $ **FLOATING
C550 vdd.n82 vss 0.02fF $ **FLOATING
C551 vdd.n83 vss 0.01fF $ **FLOATING
C552 vdd.n84 vss 0.01fF $ **FLOATING
C553 vdd.n85 vss 0.01fF $ **FLOATING
C554 vdd.n86 vss 0.01fF $ **FLOATING
C555 vdd.n87 vss 0.01fF $ **FLOATING
C556 vdd.n88 vss 0.01fF $ **FLOATING
C557 vdd.n89 vss 0.01fF $ **FLOATING
C558 vdd.n90 vss 0.01fF $ **FLOATING
C559 vdd.n91 vss 0.01fF $ **FLOATING
C560 vdd.n93 vss 0.01fF $ **FLOATING
C561 vdd.t208 vss 0.14fF
C562 vdd.t63 vss 0.14fF
C563 vdd.n94 vss 0.11fF $ **FLOATING
C564 vdd.t77 vss 0.14fF
C565 vdd.n95 vss 0.06fF $ **FLOATING
C566 vdd.t171 vss 0.14fF
C567 vdd.n96 vss 0.06fF $ **FLOATING
C568 vdd.t30 vss 0.14fF
C569 vdd.n97 vss 0.06fF $ **FLOATING
C570 vdd.t10 vss 0.14fF
C571 vdd.n98 vss 0.06fF $ **FLOATING
C572 vdd.t360 vss 0.14fF
C573 vdd.n99 vss 0.06fF $ **FLOATING
C574 vdd.t249 vss 0.14fF
C575 vdd.n100 vss 0.06fF $ **FLOATING
C576 vdd.t347 vss 0.14fF
C577 vdd.n101 vss 0.06fF $ **FLOATING
C578 vdd.t330 vss 0.14fF
C579 vdd.n102 vss 0.06fF $ **FLOATING
C580 vdd.t141 vss 0.14fF
C581 vdd.t176 vss 0.14fF
C582 vdd.n103 vss 0.11fF $ **FLOATING
C583 vdd.t195 vss 0.14fF
C584 vdd.n104 vss 0.06fF $ **FLOATING
C585 vdd.t290 vss 0.14fF
C586 vdd.n105 vss 0.06fF $ **FLOATING
C587 vdd.t307 vss 0.14fF
C588 vdd.n106 vss 0.06fF $ **FLOATING
C589 vdd.n107 vss 0.01fF $ **FLOATING
C590 vdd.n108 vss 1.31fF $ **FLOATING
C591 vdd.n109 vss 1.66fF $ **FLOATING
C592 vdd.n110 vss 0.19fF $ **FLOATING
C593 vdd.n111 vss 0.01fF $ **FLOATING
C594 vdd.n112 vss 0.42fF $ **FLOATING
C595 vdd.n113 vss 0.17fF $ **FLOATING
C596 vdd.n114 vss 0.01fF $ **FLOATING
C597 vdd.n115 vss 0.42fF $ **FLOATING
C598 vdd.n116 vss 0.16fF $ **FLOATING
C599 vdd.n117 vss 0.01fF $ **FLOATING
C600 vdd.n118 vss 0.42fF $ **FLOATING
C601 vdd.n119 vss 0.16fF $ **FLOATING
C602 vdd.n120 vss 0.01fF $ **FLOATING
C603 vdd.n121 vss 0.42fF $ **FLOATING
C604 vdd.n122 vss 0.16fF $ **FLOATING
C605 vdd.n123 vss 0.01fF $ **FLOATING
C606 vdd.n124 vss 0.42fF $ **FLOATING
C607 vdd.n125 vss 0.16fF $ **FLOATING
C608 vdd.n126 vss 0.01fF $ **FLOATING
C609 vdd.n127 vss 0.42fF $ **FLOATING
C610 vdd.n128 vss 0.16fF $ **FLOATING
C611 vdd.n129 vss 0.01fF $ **FLOATING
C612 vdd.n130 vss 0.42fF $ **FLOATING
C613 vdd.n131 vss 0.16fF $ **FLOATING
C614 vdd.n132 vss 0.01fF $ **FLOATING
C615 vdd.n133 vss 0.31fF $ **FLOATING
C616 pmos_3p3_CDNS_679510442371_1.S vss 5.22fF $ **FLOATING
C617 vdd.n134 vss 0.16fF $ **FLOATING
C618 vdd.n135 vss 0.01fF $ **FLOATING
C619 pmos_3p3_CDNS_679510442371_1.B vss 0.96fF $ **FLOATING
C620 pmos_3p3_CDNS_679510442370_1.B vss 0.97fF $ **FLOATING
C621 vdd.n136 vss 0.16fF $ **FLOATING
C622 vdd.n137 vss 0.01fF $ **FLOATING
C623 vdd.t230 vss 0.14fF
C624 vdd.t101 vss 0.14fF
C625 vdd.n138 vss 0.11fF $ **FLOATING
C626 vdd.t128 vss 0.14fF
C627 vdd.n139 vss 0.06fF $ **FLOATING
C628 vdd.t204 vss 0.14fF
C629 vdd.n140 vss 0.06fF $ **FLOATING
C630 vdd.t59 vss 0.14fF
C631 vdd.n141 vss 0.06fF $ **FLOATING
C632 vdd.t35 vss 0.14fF
C633 vdd.n142 vss 0.06fF $ **FLOATING
C634 vdd.t15 vss 0.14fF
C635 vdd.n143 vss 0.06fF $ **FLOATING
C636 vdd.t272 vss 0.14fF
C637 vdd.n144 vss 0.06fF $ **FLOATING
C638 vdd.t5 vss 0.14fF
C639 vdd.n145 vss 0.06fF $ **FLOATING
C640 vdd.t356 vss 0.14fF
C641 vdd.n146 vss 0.06fF $ **FLOATING
C642 vdd.t181 vss 0.14fF
C643 vdd.t213 vss 0.14fF
C644 vdd.n147 vss 0.11fF $ **FLOATING
C645 vdd.t221 vss 0.14fF
C646 vdd.n148 vss 0.06fF $ **FLOATING
C647 vdd.t316 vss 0.14fF
C648 vdd.n149 vss 0.06fF $ **FLOATING
C649 vdd.t339 vss 0.14fF
C650 vdd.n150 vss 0.06fF $ **FLOATING
C651 vdd.n151 vss 0.01fF $ **FLOATING
C652 vdd.n153 vss 0.01fF $ **FLOATING
C653 vdd.n154 vss 0.01fF $ **FLOATING
C654 vdd.t11 vss 1.46fF
C655 vdd.t16 vss 1.46fF
C656 vdd.t250 vss 1.46fF
C657 vdd.t6 vss 1.46fF
C658 vdd.t331 vss 1.46fF
C659 vdd.t308 vss 1.46fF
C660 vdd.t291 vss 1.46fF
C661 vdd.t196 vss 1.46fF
C662 vdd.t177 vss 1.46fF
C663 vdd.t142 vss 1.70fF
C664 vdd.n155 vss 0.01fF $ **FLOATING
C665 vdd.n157 vss 0.01fF $ **FLOATING
C666 vdd.n160 vss 0.01fF $ **FLOATING
C667 vdd.n161 vss 0.01fF $ **FLOATING
C668 vdd.n163 vss 0.01fF $ **FLOATING
C669 vdd.n165 vss 0.01fF $ **FLOATING
C670 vdd.n168 vss 0.01fF $ **FLOATING
C671 vdd.n169 vss 0.01fF $ **FLOATING
C672 vdd.n172 vss 0.01fF $ **FLOATING
C673 vdd.n173 vss 0.01fF $ **FLOATING
C674 vdd.n175 vss 0.01fF $ **FLOATING
C675 vdd.n176 vss 0.01fF $ **FLOATING
C676 vdd.n178 vss 0.01fF $ **FLOATING
C677 vdd.n179 vss 0.01fF $ **FLOATING
C678 vdd.n181 vss 0.01fF $ **FLOATING
C679 vdd.n182 vss 0.01fF $ **FLOATING
C680 vdd.n184 vss 0.01fF $ **FLOATING
C681 vdd.n185 vss 0.01fF $ **FLOATING
C682 vdd.n187 vss 0.01fF $ **FLOATING
C683 vdd.n188 vss 0.01fF $ **FLOATING
C684 vdd.n189 vss 0.01fF $ **FLOATING
C685 vdd.n191 vss 0.01fF $ **FLOATING
C686 vdd.n192 vss 0.01fF $ **FLOATING
C687 vdd.n193 vss 0.01fF $ **FLOATING
C688 vdd.n194 vss 0.01fF $ **FLOATING
C689 vdd.n195 vss 0.01fF $ **FLOATING
C690 vdd.n196 vss 0.01fF $ **FLOATING
C691 vdd.n197 vss 0.01fF $ **FLOATING
C692 vdd.n198 vss 0.01fF $ **FLOATING
C693 vdd.n199 vss 0.01fF $ **FLOATING
C694 vdd.n200 vss 0.01fF $ **FLOATING
C695 vdd.n201 vss 0.01fF $ **FLOATING
C696 vdd.n202 vss 0.01fF $ **FLOATING
C697 vdd.n203 vss 0.01fF $ **FLOATING
C698 vdd.n204 vss 0.31fF $ **FLOATING
C699 vdd.n206 vss 0.31fF $ **FLOATING
C700 vdd.n207 vss 0.01fF $ **FLOATING
C701 vdd.n208 vss 0.01fF $ **FLOATING
C702 vdd.n209 vss 0.01fF $ **FLOATING
C703 vdd.n210 vss 0.01fF $ **FLOATING
C704 vdd.n211 vss 0.01fF $ **FLOATING
C705 vdd.n212 vss 0.01fF $ **FLOATING
C706 vdd.n213 vss 0.01fF $ **FLOATING
C707 vdd.n214 vss 0.01fF $ **FLOATING
C708 vdd.n215 vss 0.01fF $ **FLOATING
C709 vdd.n216 vss 0.01fF $ **FLOATING
C710 vdd.n217 vss 0.38fF $ **FLOATING
C711 vdd.n218 vss 0.02fF $ **FLOATING
C712 vdd.n219 vss 1.05fF $ **FLOATING
C713 vdd.n221 vss 0.01fF $ **FLOATING
C714 vdd.n222 vss 0.01fF $ **FLOATING
C715 vdd.n223 vss 0.02fF $ **FLOATING
C716 vdd.n224 vss 0.02fF $ **FLOATING
C717 vdd.n225 vss 0.20fF $ **FLOATING
C718 vdd.n226 vss 0.20fF $ **FLOATING
C719 vdd.n227 vss 0.22fF $ **FLOATING
C720 vdd.t286 vss 1.46fF
C721 vdd.t26 vss 1.46fF
C722 vdd.t40 vss 1.46fF
C723 vdd.t321 vss 1.46fF
C724 vdd.t55 vss 1.46fF
C725 vdd.t88 vss 1.46fF
C726 vdd.t120 vss 1.62fF
C727 vdd.n228 vss 0.97fF $ **FLOATING
C728 vdd.n229 vss 0.21fF $ **FLOATING
C729 vdd.n230 vss 0.21fF $ **FLOATING
C730 vdd.n231 vss 0.05fF $ **FLOATING
C731 vdd.n232 vss 1.23fF $ **FLOATING
C732 vdd.n233 vss 0.93fF $ **FLOATING
C733 vdd.n234 vss 0.48fF $ **FLOATING
C734 vdd.n235 vss 0.18fF $ **FLOATING
C735 vdd.n236 vss 0.01fF $ **FLOATING
C736 vdd.n237 vss 0.42fF $ **FLOATING
C737 vdd.n238 vss 0.17fF $ **FLOATING
C738 vdd.n239 vss 0.01fF $ **FLOATING
C739 vdd.n240 vss 0.42fF $ **FLOATING
C740 vdd.n241 vss 0.16fF $ **FLOATING
C741 vdd.n242 vss 0.01fF $ **FLOATING
C742 vdd.n243 vss 0.42fF $ **FLOATING
C743 vdd.n244 vss 0.16fF $ **FLOATING
C744 vdd.n245 vss 0.01fF $ **FLOATING
C745 vdd.n246 vss 0.42fF $ **FLOATING
C746 vdd.n247 vss 0.16fF $ **FLOATING
C747 vdd.n248 vss 0.01fF $ **FLOATING
C748 vdd.n249 vss 0.42fF $ **FLOATING
C749 vdd.n250 vss 0.16fF $ **FLOATING
C750 vdd.n251 vss 0.01fF $ **FLOATING
C751 vdd.n252 vss 0.42fF $ **FLOATING
C752 vdd.n253 vss 0.16fF $ **FLOATING
C753 vdd.n254 vss 0.01fF $ **FLOATING
C754 vdd.n255 vss 0.42fF $ **FLOATING
C755 vdd.n256 vss 0.42fF $ **FLOATING
C756 pmos_3p3_CDNS_679510442370_1.S vss 5.49fF $ **FLOATING
C757 vdd.n257 vss 0.16fF $ **FLOATING
C758 vdd.n258 vss 0.01fF $ **FLOATING
C759 vdd.n259 vss 0.16fF $ **FLOATING
C760 vdd.n260 vss 0.01fF $ **FLOATING
C761 vdd.n261 vss 0.16fF $ **FLOATING
C762 vdd.n262 vss 0.01fF $ **FLOATING
C763 vdd.n263 vss 0.42fF $ **FLOATING
C764 vdd.n264 vss 0.16fF $ **FLOATING
C765 vdd.n265 vss 0.01fF $ **FLOATING
C766 vdd.n266 vss 0.42fF $ **FLOATING
C767 vdd.n267 vss 0.16fF $ **FLOATING
C768 vdd.n268 vss 0.01fF $ **FLOATING
C769 vdd.n269 vss 0.42fF $ **FLOATING
C770 vdd.n270 vss 0.16fF $ **FLOATING
C771 vdd.n271 vss 0.01fF $ **FLOATING
C772 vdd.n272 vss 0.42fF $ **FLOATING
C773 vdd.n273 vss 0.16fF $ **FLOATING
C774 vdd.n274 vss 0.01fF $ **FLOATING
C775 vdd.n275 vss 0.42fF $ **FLOATING
C776 vdd.n276 vss 0.16fF $ **FLOATING
C777 vdd.n277 vss 0.01fF $ **FLOATING
C778 vdd.n278 vss 0.42fF $ **FLOATING
C779 vdd.n279 vss 0.16fF $ **FLOATING
C780 vdd.n280 vss 0.01fF $ **FLOATING
C781 vdd.n281 vss 0.42fF $ **FLOATING
C782 vdd.n282 vss 0.16fF $ **FLOATING
C783 vdd.n283 vss 0.01fF $ **FLOATING
C784 vdd.n284 vss 0.42fF $ **FLOATING
C785 vdd.n285 vss 0.42fF $ **FLOATING
C786 vdd.n286 vss 0.33fF $ **FLOATING
C787 vdd.n287 vss 0.01fF $ **FLOATING
C788 vdd.n288 vss 0.16fF $ **FLOATING
C789 vdd.n289 vss 0.17fF $ **FLOATING
C790 vdd.t31 vss 1.46fF
C791 vdd.t172 vss 1.46fF
C792 vdd.t78 vss 1.46fF
C793 vdd.t64 vss 1.46fF
C794 vdd.t209 vss 1.34fF
C795 vdd.n290 vss 0.92fF $ **FLOATING
C796 vdd.n291 vss 0.14fF $ **FLOATING
C797 vdd.n292 vss 0.01fF $ **FLOATING
C798 vdd.n293 vss 0.42fF $ **FLOATING
C799 vdd.n294 vss 0.16fF $ **FLOATING
C800 vdd.n295 vss 0.01fF $ **FLOATING
C801 vdd.n296 vss 0.42fF $ **FLOATING
C802 vdd.n297 vss 0.16fF $ **FLOATING
C803 vdd.n298 vss 0.01fF $ **FLOATING
C804 vdd.n299 vss 0.42fF $ **FLOATING
C805 vdd.n300 vss 0.16fF $ **FLOATING
C806 vdd.n301 vss 0.01fF $ **FLOATING
C807 vdd.n302 vss 0.42fF $ **FLOATING
C808 vdd.n303 vss 0.16fF $ **FLOATING
C809 vdd.n304 vss 0.01fF $ **FLOATING
C810 vdd.n305 vss 0.42fF $ **FLOATING
C811 vdd.n306 vss 0.16fF $ **FLOATING
C812 vdd.n307 vss 0.01fF $ **FLOATING
C813 vdd.n308 vss 0.42fF $ **FLOATING
C814 vdd.n309 vss 0.16fF $ **FLOATING
C815 vdd.n310 vss 0.01fF $ **FLOATING
C816 vdd.n311 vss 0.42fF $ **FLOATING
C817 vdd.n312 vss 0.16fF $ **FLOATING
C818 vdd.n313 vss 0.01fF $ **FLOATING
C819 vdd.n314 vss 0.42fF $ **FLOATING
C820 vdd.n315 vss 0.42fF $ **FLOATING
C821 vdd.n316 vss 0.16fF $ **FLOATING
C822 vdd.n317 vss 0.01fF $ **FLOATING
C823 vdd.n318 vss 0.16fF $ **FLOATING
C824 vdd.n319 vss 0.01fF $ **FLOATING
C825 vdd.n320 vss 0.17fF $ **FLOATING
C826 vdd.n321 vss 0.42fF $ **FLOATING
C827 vdd.n322 vss 0.08fF $ **FLOATING
C828 vdd.n323 vss 0.08fF $ **FLOATING
C829 vdd.n324 vss 0.08fF $ **FLOATING
C830 vdd.n325 vss 0.08fF $ **FLOATING
C831 vdd.n326 vss 0.07fF $ **FLOATING
C832 vdd.n327 vss 0.08fF $ **FLOATING
C833 vdd.n328 vss 0.08fF $ **FLOATING
C834 vdd.n329 vss 0.09fF $ **FLOATING
C835 vdd.n330 vss 0.01fF $ **FLOATING
C836 vdd.n331 vss 0.01fF $ **FLOATING
C837 vdd.n332 vss 0.01fF $ **FLOATING
C838 vdd.n333 vss 0.01fF $ **FLOATING
C839 vdd.n334 vss 0.01fF $ **FLOATING
C840 vdd.n335 vss 0.01fF $ **FLOATING
C841 vdd.n336 vss 0.01fF $ **FLOATING
C842 vdd.n338 vss 0.01fF $ **FLOATING
C843 vdd.n339 vss 0.01fF $ **FLOATING
C844 vdd.n340 vss 0.01fF $ **FLOATING
C845 vdd.n341 vss 2.69fF $ **FLOATING
C846 vdd.t557 vss 5.04fF
C847 vdd.t368 vss 6.46fF
C848 vdd.t560 vss 7.35fF
C849 vdd.t558 vss 7.35fF
C850 vdd.t559 vss 6.26fF
C851 vdd.t378 vss 6.26fF
C852 vdd.t410 vss 6.26fF
C853 vdd.t372 vss 6.26fF
C854 vdd.t369 vss 6.26fF
C855 vdd.t400 vss 5.00fF
C856 vdd.n342 vss 2.71fF $ **FLOATING
C857 vdd.n343 vss 1.86fF $ **FLOATING
C858 vdd.n344 vss 8.91fF $ **FLOATING
C859 vdd.t375 vss 3.23fF
C860 vdd.n345 vss 1.26fF $ **FLOATING
C861 vdd.n346 vss 0.07fF $ **FLOATING
C862 vdd.n347 vss 0.76fF $ **FLOATING
C863 vdd.t407 vss 3.45fF
C864 vdd.n348 vss 3.13fF $ **FLOATING
C865 vdd.n349 vss 0.13fF $ **FLOATING
C866 vdd.n350 vss 2.10fF $ **FLOATING
C867 vdd.t392 vss 4.09fF
C868 vdd.n351 vss 1.80fF $ **FLOATING
C869 vdd.n352 vss 0.09fF $ **FLOATING
C870 vdd.n353 vss 1.48fF $ **FLOATING
C871 vdd.n354 vss 0.27fF $ **FLOATING
C872 vdd.n355 vss 1.67fF $ **FLOATING
C873 vdd.n356 vss 0.03fF $ **FLOATING
C874 vdd.n357 vss 0.31fF $ **FLOATING
C875 vdd.n358 vss 2.79fF $ **FLOATING
C876 vdd.n359 vss 0.05fF $ **FLOATING
C877 vdd.t50 vss 8.34fF
C878 vdd.t69 vss 8.34fF
C879 vdd.t110 vss 6.13fF
C880 vdd.n360 vss 4.17fF $ **FLOATING
C881 vdd.n361 vss 0.45fF $ **FLOATING
C882 vdd.t137 vss 2.58fF
C883 vdd.t594 vss 0.23fF
C884 vdd.t561 vss 2.24fF
C885 vdd.t83 vss 4.11fF
C886 vdd.t255 vss 1.99fF
C887 vdd.t186 vss 0.48fF
C888 vdd.t115 vss 1.87fF
C889 vdd.t254 vss 0.22fF
C890 vdd.t82 vss 0.10fF
C891 vdd.t92 vss 0.10fF
C892 vdd.t136 vss 0.11fF
C893 vdd.t150 vss 0.11fF
C894 vdd.n362 vss 0.13fF $ **FLOATING
C895 vdd.n363 vss 0.17fF $ **FLOATING
C896 vdd.t185 vss 0.22fF
C897 vdd.t163 vss 0.10fF
C898 vdd.t217 vss 0.10fF
C899 vdd.t259 vss 0.10fF
C900 vdd.t299 vss 0.10fF
C901 vdd.t0 vss 0.30fF
C902 vdd.t146 vss 0.30fF
C903 vdd.t73 vss 0.30fF
C904 vdd.t105 vss 0.30fF
C905 vdd.t132 vss 0.30fF
C906 vdd.t159 vss 0.30fF
C907 vdd.t364 vss 0.50fF
C908 vdd.t200 vss 0.64fF
C909 vdd.n364 vss 0.24fF $ **FLOATING
C910 vdd.n365 vss 0.24fF $ **FLOATING
C911 vdd.n366 vss 0.24fF $ **FLOATING
C912 vdd.n367 vss 0.24fF $ **FLOATING
C913 vdd.n368 vss 0.24fF $ **FLOATING
C914 vdd.n369 vss 0.23fF $ **FLOATING
C915 vdd.n370 vss 0.11fF $ **FLOATING
C916 vdd.n371 vss 0.10fF $ **FLOATING
C917 vdd.n372 vss 0.10fF $ **FLOATING
C918 vdd.n373 vss 0.11fF $ **FLOATING
C919 vdd.t343 vss 0.15fF
C920 vdd.n374 vss 0.38fF $ **FLOATING
C921 vdd.t268 vss 0.18fF
C922 vdd.t114 vss 0.21fF
C923 vdd.t295 vss 0.15fF
C924 vdd.n375 vss 0.13fF $ **FLOATING
C925 vdd.t276 vss 0.13fF
C926 vdd.n376 vss 0.37fF $ **FLOATING
C927 vdd.t303 vss 0.08fF
C928 vdd.t124 vss 0.10fF
C929 vdd.t167 vss 0.10fF
C930 vdd.t239 vss 0.10fF
C931 vdd.t263 vss 0.10fF
C932 vdd.t335 vss 0.30fF
C933 vdd.t96 vss 0.30fF
C934 vdd.t20 vss 0.30fF
C935 vdd.t49 vss 0.30fF
C936 vdd.t68 vss 0.30fF
C937 vdd.t109 vss 0.30fF
C938 vdd.t312 vss 0.50fF
C939 vdd.t154 vss 0.64fF
C940 vdd.n377 vss 0.24fF $ **FLOATING
C941 vdd.n378 vss 0.24fF $ **FLOATING
C942 vdd.n379 vss 0.24fF $ **FLOATING
C943 vdd.n380 vss 0.24fF $ **FLOATING
C944 vdd.n381 vss 0.24fF $ **FLOATING
C945 vdd.n382 vss 0.23fF $ **FLOATING
C946 vdd.n383 vss 0.11fF $ **FLOATING
C947 vdd.n384 vss 0.10fF $ **FLOATING
C948 vdd.n385 vss 0.10fF $ **FLOATING
C949 vdd.n386 vss 0.10fF $ **FLOATING
C950 vdd.n387 vss 0.08fF $ **FLOATING
C951 vdd.n388 vss 0.35fF $ **FLOATING
C952 vdd.n389 vss 29.01fF $ **FLOATING
C953 vdd.t21 vss 8.34fF
C954 vdd.t97 vss 8.34fF
C955 vdd.t1 vss 6.17fF
C956 vdd.t240 vss 3.94fF
C957 vdd.t453 vss 1.59fF
C958 vdd.t494 vss 0.88fF
C959 vdd.t264 vss 2.11fF
C960 vdd.n390 vss 3.29fF $ **FLOATING
C961 vdd.n391 vss 0.83fF $ **FLOATING
C962 vdd.n392 vss 0.22fF $ **FLOATING
C963 vdd.n393 vss 6.87fF $ **FLOATING
C964 vdd.n394 vss 0.45fF $ **FLOATING
C965 vdd.t539 vss 1.09fF
C966 vdd.t547 vss 1.90fF
C967 vdd.n395 vss 3.96fF $ **FLOATING
C968 vdd.t155 vss 2.36fF
C969 vdd.n396 vss 2.08fF $ **FLOATING
C970 vdd.n397 vss 0.21fF $ **FLOATING
C971 vdd.n398 vss 0.21fF $ **FLOATING
C972 vdd.t527 vss 1.46fF
C973 vdd.t524 vss 1.46fF
C974 vdd.t521 vss 1.46fF
C975 vdd.t554 vss 1.46fF
C976 vdd.t529 vss 1.46fF
C977 vdd.t553 vss 1.46fF
C978 vdd.t551 vss 2.30fF
C979 vdd.t538 vss 0.85fF
C980 vdd.n399 vss 0.83fF $ **FLOATING
C981 vdd.t549 vss 1.06fF
C982 vdd.t542 vss 1.46fF
C983 vdd.t552 vss 1.46fF
C984 vdd.t555 vss 1.46fF
C985 vdd.t522 vss 1.46fF
C986 vdd.t520 vss 1.46fF
C987 vdd.t523 vss 0.97fF
C988 vdd.n400 vss 1.81fF $ **FLOATING
C989 vdd.n401 vss 0.38fF $ **FLOATING
C990 vdd.n402 vss 0.38fF $ **FLOATING
C991 vdd.t545 vss 1.46fF
C992 vdd.t506 vss 1.46fF
C993 vdd.t531 vss 2.54fF
C994 vdd.t544 vss 2.54fF
C995 vdd.t550 vss 1.46fF
C996 vdd.t540 vss 1.46fF
C997 vdd.t536 vss 1.46fF
C998 vdd.t534 vss 1.46fF
C999 vdd.t526 vss 1.06fF
C1000 vdd.t505 vss 1.46fF
C1001 vdd.t537 vss 1.46fF
C1002 vdd.t528 vss 2.54fF
C1003 vdd.t556 vss 2.54fF
C1004 vdd.t530 vss 1.46fF
C1005 vdd.t532 vss 1.46fF
C1006 vdd.t533 vss 1.13fF
C1007 vdd.n403 vss 0.73fF $ **FLOATING
C1008 vdd.n404 vss 0.45fF $ **FLOATING
C1009 vdd.n405 vss 0.45fF $ **FLOATING
C1010 vdd.t397 vss 2.40fF
C1011 vdd.t535 vss 1.46fF
C1012 vdd.t541 vss 1.46fF
C1013 vdd.t543 vss 1.46fF
C1014 vdd.t546 vss 1.46fF
C1015 vdd.t519 vss 1.46fF
C1016 vdd.t548 vss 1.46fF
C1017 vdd.t525 vss 3.30fF
C1018 vdd.n406 vss 3.02fF $ **FLOATING
C1019 vdd.n407 vss 0.29fF $ **FLOATING
C1020 vdd.n408 vss 0.30fF $ **FLOATING
C1021 vdd.n409 vss 1.53fF $ **FLOATING
C1022 vdd.t383 vss 0.84fF
C1023 vdd.n410 vss 1.18fF $ **FLOATING
C1024 vdd.n411 vss 0.03fF $ **FLOATING
C1025 vdd.n412 vss 0.31fF $ **FLOATING
C1026 vdd.n413 vss 1.33fF $ **FLOATING
C1027 vdd.n414 vss 0.03fF $ **FLOATING
C1028 vdd.n415 vss 0.31fF $ **FLOATING
C1029 vdd.n417 vss 26.84fF $ **FLOATING
C1030 vdd.n418 vss 27.56fF $ **FLOATING
C1031 vdd.n420 vss 1.45fF $ **FLOATING
C1032 vdd.n422 vss 0.32fF $ **FLOATING
C1033 vdd.n423 vss 0.47fF $ **FLOATING
C1034 vdd.n425 vss 0.37fF $ **FLOATING
C1035 vdd.n427 vss 0.39fF $ **FLOATING
C1036 vdd.n429 vss 0.37fF $ **FLOATING
C1037 vdd.n431 vss 0.37fF $ **FLOATING
C1038 vdd.n433 vss 0.38fF $ **FLOATING
C1039 vdd.n434 vss 0.38fF $ **FLOATING
C1040 vdd.n437 vss 0.36fF $ **FLOATING
C1041 vdd.n439 vss 0.30fF $ **FLOATING
C1042 vdd.n441 vss 0.34fF $ **FLOATING
C1043 vdd.n443 vss 0.34fF $ **FLOATING
C1044 vdd.n444 vss 0.52fF $ **FLOATING
C1045 vdd.n446 vss 0.34fF $ **FLOATING
C1046 vdd.n448 vss 20.49fF $ **FLOATING
C1047 vdd.n449 vss 20.47fF $ **FLOATING
C1048 vdd.n451 vss 0.28fF $ **FLOATING
C1049 vdd.n453 vss 0.30fF $ **FLOATING
C1050 vdd.n454 vss 0.30fF $ **FLOATING
C1051 vdd.n456 vss 0.30fF $ **FLOATING
C1052 vdd.n458 vss 0.36fF $ **FLOATING
C1053 vdd.n460 vss 45.02fF $ **FLOATING
C1054 vdd.n461 vss 45.02fF $ **FLOATING
C1055 vdd.n463 vss 0.37fF $ **FLOATING
C1056 vdd.n465 vss 0.28fF $ **FLOATING
C1057 vdd.n467 vss 0.30fF $ **FLOATING
C1058 vdd.n469 vss 0.30fF $ **FLOATING
C1059 vdd.n471 vss 0.39fF $ **FLOATING
C1060 vdd.n473 vss 0.30fF $ **FLOATING
C1061 vdd.n475 vss 6.26fF $ **FLOATING
C1062 vdd.n476 vss 0.02fF $ **FLOATING
C1063 vdd.n477 vss 0.00fF $ **FLOATING
C1064 vdd.n478 vss 0.02fF $ **FLOATING
C1065 vdd.n479 vss 3.66fF $ **FLOATING
C1066 vdd.n480 vss 0.18fF $ **FLOATING
C1067 vdd.n481 vss 0.00fF $ **FLOATING
C1068 vdd.n482 vss 0.01fF $ **FLOATING
C1069 vdd.n483 vss 0.00fF $ **FLOATING
C1070 vdd.n484 vss 0.02fF $ **FLOATING
C1071 vdd.n485 vss 0.88fF $ **FLOATING
C1072 vdd.n486 vss 1.54fF $ **FLOATING
C1073 vdd.n487 vss 1.60fF $ **FLOATING
C1074 vdd.n488 vss 0.00fF $ **FLOATING
C1075 vdd.n489 vss 0.10fF $ **FLOATING
C1076 vdd.n490 vss 0.01fF $ **FLOATING
C1077 vdd.n491 vss 0.02fF $ **FLOATING
C1078 vdd.n492 vss 0.02fF $ **FLOATING
C1079 vdd.n493 vss 0.17fF $ **FLOATING
C1080 vdd.n494 vss 0.03fF $ **FLOATING
C1081 vdd.n495 vss 0.01fF $ **FLOATING
C1082 vdd.n496 vss 0.04fF $ **FLOATING
C1083 vdd.n497 vss 0.02fF $ **FLOATING
C1084 vdd.n498 vss 1.64fF $ **FLOATING
C1085 vdd.n499 vss 0.25fF $ **FLOATING
C1086 vdd.n500 vss 1.40fF $ **FLOATING
C1087 vdd.n502 vss 10.58fF $ **FLOATING
C1088 vdd.n503 vss 8.28fF $ **FLOATING
C1089 vdd.n505 vss 3.09fF $ **FLOATING
C1090 vdd.n506 vss 0.80fF $ **FLOATING
C1091 vdd.n507 vss 0.02fF $ **FLOATING
C1092 vdd.n508 vss 0.02fF $ **FLOATING
C1093 vdd.n510 vss 1.82fF $ **FLOATING
C1094 vdd.n511 vss 1.82fF $ **FLOATING
C1095 vdd.n512 vss 3.09fF $ **FLOATING
C1096 vdd.n513 vss 0.80fF $ **FLOATING
C1097 vdd.n514 vss 0.02fF $ **FLOATING
C1098 vdd.n515 vss 0.02fF $ **FLOATING
C1099 vdd.n517 vss 5.55fF $ **FLOATING
C1100 vdd.n518 vss 5.56fF $ **FLOATING
C1101 vdd.n519 vss 0.02fF $ **FLOATING
C1102 vdd.n520 vss 0.00fF $ **FLOATING
C1103 vdd.n521 vss 0.01fF $ **FLOATING
C1104 vdd.n522 vss 0.01fF $ **FLOATING
C1105 vdd.n523 vss 3.63fF $ **FLOATING
C1106 vdd.n524 vss 0.21fF $ **FLOATING
C1107 vdd.n526 vss 0.01fF $ **FLOATING
C1108 vdd.n528 vss 1.86fF $ **FLOATING
C1109 vdd.n529 vss 1.86fF $ **FLOATING
C1110 vdd.n531 vss 0.01fF $ **FLOATING
C1111 vdd.n533 vss 4.41fF $ **FLOATING
C1112 vdd.n534 vss 4.41fF $ **FLOATING
C1113 vdd.n536 vss 0.02fF $ **FLOATING
C1114 vdd.n538 vss 2.00fF $ **FLOATING
C1115 vdd.n539 vss 2.08fF $ **FLOATING
C1116 vdd.n541 vss 0.23fF $ **FLOATING
C1117 vdd.n542 vss 0.39fF $ **FLOATING
C1118 vdd.n543 vss 6.26fF $ **FLOATING
C1119 vdd.n545 vss 14.62fF $ **FLOATING
C1120 vdd.n546 vss 14.64fF $ **FLOATING
C1121 vdd.n548 vss 0.34fF $ **FLOATING
C1122 vdd.n550 vss 0.34fF $ **FLOATING
C1123 vdd.n551 vss 0.34fF $ **FLOATING
C1124 vdd.n553 vss 3.01fF $ **FLOATING
C1125 vdd.n554 vss 15.63fF $ **FLOATING
C1126 vdd.n556 vss 0.34fF $ **FLOATING
C1127 vdd.n558 vss 0.34fF $ **FLOATING
C1128 vdd.n560 vss 0.34fF $ **FLOATING
C1129 vdd.n562 vss 0.34fF $ **FLOATING
C1130 vdd.n564 vss 0.34fF $ **FLOATING
C1131 vdd.n566 vss 0.34fF $ **FLOATING
C1132 vdd.n568 vss 0.34fF $ **FLOATING
C1133 vdd.n570 vss 0.34fF $ **FLOATING
C1134 vdd.n572 vss 0.34fF $ **FLOATING
C1135 vdd.n574 vss 0.34fF $ **FLOATING
C1136 vdd.n576 vss 0.34fF $ **FLOATING
C1137 vdd.n577 vss 12.14fF $ **FLOATING
C1138 vdd.n579 vss 1.37fF $ **FLOATING
C1139 vdd.n581 vss 33.51fF $ **FLOATING
C1140 vdd.n582 vss 46.89fF $ **FLOATING
C1141 vdd.n583 vss 3.81fF $ **FLOATING
C1142 vdd.t511 vss 2.67fF
C1143 vdd.t516 vss 0.46fF
C1144 vdd.t518 vss 0.46fF
C1145 vdd.t513 vss 0.46fF
C1146 vdd.t515 vss 0.46fF
C1147 vdd.t508 vss 0.46fF
C1148 vdd.t512 vss 0.46fF
C1149 vdd.t517 vss 0.46fF
C1150 vdd.t510 vss 0.37fF
C1151 vdd.n584 vss 0.93fF $ **FLOATING
C1152 vdd.n585 vss 0.23fF $ **FLOATING
C1153 vdd.t514 vss 0.15fF
C1154 vdd.n586 vss 0.19fF $ **FLOATING
C1155 vdd.n587 vss 0.52fF $ **FLOATING
C1156 vdd.n588 vss 0.50fF $ **FLOATING
C1157 vdd.n589 vss 0.18fF $ **FLOATING
C1158 vdd.t507 vss 0.27fF
C1159 vdd.n590 vss 1.05fF $ **FLOATING
C1160 vdd.n591 vss 0.97fF $ **FLOATING
C1161 vdd.n592 vss 2.63fF $ **FLOATING
C1162 vdd.t630 vss 0.01fF
C1163 vdd.t601 vss 0.01fF
C1164 vdd.t638 vss 0.01fF
C1165 vdd.t623 vss 0.01fF
C1166 vdd.t667 vss 0.01fF
C1167 vdd.t642 vss 0.02fF
C1168 vdd.n593 vss 0.04fF $ **FLOATING
C1169 vdd.n594 vss 0.03fF $ **FLOATING
C1170 vdd.n595 vss 0.03fF $ **FLOATING
C1171 vdd.n596 vss 0.03fF $ **FLOATING
C1172 vdd.n597 vss 0.02fF $ **FLOATING
C1173 vdd.t648 vss 0.01fF
C1174 vdd.t609 vss 0.01fF
C1175 vdd.t628 vss 0.01fF
C1176 vdd.t682 vss 0.01fF
C1177 vdd.t606 vss 0.01fF
C1178 vdd.t633 vss 0.02fF
C1179 vdd.n598 vss 0.04fF $ **FLOATING
C1180 vdd.n599 vss 0.03fF $ **FLOATING
C1181 vdd.n600 vss 0.03fF $ **FLOATING
C1182 vdd.n601 vss 0.03fF $ **FLOATING
C1183 vdd.n602 vss 0.02fF $ **FLOATING
C1184 vdd.n603 vss 0.01fF $ **FLOATING
C1185 vin2.t69 vss 0.30fF
C1186 vin2.t18 vss 0.30fF
C1187 vin2.t79 vss 0.30fF
C1188 vin2.t23 vss 0.30fF
C1189 vin2.t28 vss 0.30fF
C1190 vin2.t30 vss 0.30fF
C1191 vin2.t39 vss 0.30fF
C1192 vin2.t24 vss 0.30fF
C1193 vin2.t48 vss 0.30fF
C1194 vin2.t52 vss 0.30fF
C1195 vin2.t76 vss 0.28fF
C1196 vin2.t72 vss 0.28fF
C1197 vin2.t67 vss 0.28fF
C1198 vin2.t42 vss 0.28fF
C1199 vin2.t35 vss 0.28fF
C1200 vin2.t60 vss 0.28fF
C1201 vin2.t0 vss 0.28fF
C1202 vin2.t55 vss 0.28fF
C1203 vin2.t50 vss 0.28fF
C1204 vin2.t47 vss 0.28fF
C1205 vin2.t68 vss 0.28fF
C1206 vin2.t44 vss 0.28fF
C1207 vin2.t36 vss 0.28fF
C1208 vin2.t31 vss 0.28fF
C1209 vin2.t11 vss 0.28fF
C1210 vin2.t25 vss 0.29fF
C1211 vin2.n0 vss 0.27fF $ **FLOATING
C1212 vin2.n1 vss 0.15fF $ **FLOATING
C1213 vin2.n2 vss 0.15fF $ **FLOATING
C1214 vin2.n3 vss 0.15fF $ **FLOATING
C1215 vin2.n4 vss 0.15fF $ **FLOATING
C1216 vin2.n5 vss 0.15fF $ **FLOATING
C1217 vin2.n6 vss 0.15fF $ **FLOATING
C1218 vin2.n7 vss 0.15fF $ **FLOATING
C1219 vin2.n8 vss 0.19fF $ **FLOATING
C1220 vin2.n9 vss 0.19fF $ **FLOATING
C1221 vin2.n10 vss 0.15fF $ **FLOATING
C1222 vin2.n11 vss 0.15fF $ **FLOATING
C1223 vin2.n12 vss 0.15fF $ **FLOATING
C1224 vin2.n13 vss 0.15fF $ **FLOATING
C1225 vin2.n14 vss 0.14fF $ **FLOATING
C1226 vin2.t3 vss 0.28fF
C1227 vin2.t59 vss 0.28fF
C1228 vin2.t7 vss 0.28fF
C1229 vin2.t10 vss 0.29fF
C1230 vin2.n15 vss 0.27fF $ **FLOATING
C1231 vin2.n16 vss 0.15fF $ **FLOATING
C1232 vin2.n17 vss 0.14fF $ **FLOATING
C1233 vin2.n18 vss 0.61fF $ **FLOATING
C1234 vin2.t73 vss 0.30fF
C1235 vin2.t77 vss 0.30fF
C1236 vin2.t75 vss 0.30fF
C1237 vin2.t1 vss 0.30fF
C1238 vin2.t8 vss 0.30fF
C1239 vin2.t29 vss 0.30fF
C1240 vin2.t15 vss 0.30fF
C1241 vin2.t34 vss 0.30fF
C1242 vin2.t32 vss 0.30fF
C1243 vin2.t21 vss 0.31fF
C1244 vin2.n19 vss 0.32fF $ **FLOATING
C1245 vin2.n20 vss 0.17fF $ **FLOATING
C1246 vin2.n21 vss 0.17fF $ **FLOATING
C1247 vin2.n22 vss 0.17fF $ **FLOATING
C1248 vin2.n23 vss 0.17fF $ **FLOATING
C1249 vin2.n24 vss 0.17fF $ **FLOATING
C1250 vin2.n25 vss 0.17fF $ **FLOATING
C1251 vin2.n26 vss 0.17fF $ **FLOATING
C1252 vin2.n27 vss 0.29fF $ **FLOATING
C1253 vin2.n28 vss 1.21fF $ **FLOATING
C1254 vin2.n29 vss 0.62fF $ **FLOATING
C1255 vin2.n30 vss 0.17fF $ **FLOATING
C1256 vin2.n31 vss 0.17fF $ **FLOATING
C1257 vin2.n32 vss 0.17fF $ **FLOATING
C1258 vin2.n33 vss 0.17fF $ **FLOATING
C1259 vin2.n34 vss 0.17fF $ **FLOATING
C1260 vin2.n35 vss 0.17fF $ **FLOATING
C1261 vin2.n36 vss 0.17fF $ **FLOATING
C1262 vin2.n37 vss 0.17fF $ **FLOATING
C1263 vin2.n38 vss 0.55fF $ **FLOATING
C1264 vin2.t71 vss 0.28fF
C1265 vin2.t13 vss 0.28fF
C1266 vin2.t37 vss 0.28fF
C1267 vin2.t9 vss 0.28fF
C1268 vin2.t26 vss 0.28fF
C1269 vin2.t56 vss 0.28fF
C1270 vin2.t65 vss 0.28fF
C1271 vin2.t16 vss 0.28fF
C1272 vin2.t62 vss 0.28fF
C1273 vin2.t4 vss 0.30fF
C1274 vin2.n39 vss 0.26fF $ **FLOATING
C1275 vin2.n40 vss 0.14fF $ **FLOATING
C1276 vin2.n41 vss 0.14fF $ **FLOATING
C1277 vin2.n42 vss 0.14fF $ **FLOATING
C1278 vin2.n43 vss 0.14fF $ **FLOATING
C1279 vin2.n44 vss 0.14fF $ **FLOATING
C1280 vin2.n45 vss 0.14fF $ **FLOATING
C1281 vin2.n46 vss 0.14fF $ **FLOATING
C1282 vin2.n47 vss 0.47fF $ **FLOATING
C1283 vin2.t43 vss 0.28fF
C1284 vin2.t19 vss 0.28fF
C1285 vin2.t58 vss 0.28fF
C1286 vin2.t33 vss 0.28fF
C1287 vin2.t12 vss 0.28fF
C1288 vin2.t41 vss 0.28fF
C1289 vin2.t40 vss 0.28fF
C1290 vin2.t74 vss 0.28fF
C1291 vin2.t54 vss 0.28fF
C1292 vin2.t2 vss 0.30fF
C1293 vin2.n48 vss 0.26fF $ **FLOATING
C1294 vin2.n49 vss 0.14fF $ **FLOATING
C1295 vin2.n50 vss 0.14fF $ **FLOATING
C1296 vin2.n51 vss 0.14fF $ **FLOATING
C1297 vin2.n52 vss 0.14fF $ **FLOATING
C1298 vin2.n53 vss 0.14fF $ **FLOATING
C1299 vin2.n54 vss 0.14fF $ **FLOATING
C1300 vin2.n55 vss 0.14fF $ **FLOATING
C1301 vin2.n56 vss 0.19fF $ **FLOATING
C1302 vin2.n57 vss 4.30fF $ **FLOATING
C1303 vin2.t53 vss 0.28fF
C1304 vin2.t46 vss 0.28fF
C1305 vin2.t14 vss 0.28fF
C1306 vin2.t38 vss 0.28fF
C1307 vin2.t61 vss 0.28fF
C1308 vin2.t27 vss 0.28fF
C1309 vin2.t57 vss 0.28fF
C1310 vin2.t66 vss 0.28fF
C1311 vin2.t17 vss 0.28fF
C1312 vin2.t63 vss 0.28fF
C1313 vin2.n58 vss 0.01fF $ **FLOATING
C1314 vin2.n59 vss 0.01fF $ **FLOATING
C1315 vin2.t64 vss 0.28fF
C1316 vin2.t5 vss 0.28fF
C1317 vin2.t49 vss 0.28fF
C1318 vin2.t78 vss 0.28fF
C1319 vin2.t20 vss 0.28fF
C1320 vin2.t45 vss 0.28fF
C1321 vin2.t6 vss 0.28fF
C1322 vin2.t22 vss 0.28fF
C1323 vin2.t51 vss 0.28fF
C1324 vin2.t70 vss 0.30fF
C1325 vin2.n60 vss 0.26fF $ **FLOATING
C1326 vin2.n61 vss 0.14fF $ **FLOATING
C1327 vin2.n62 vss 0.14fF $ **FLOATING
C1328 vin2.n63 vss 0.14fF $ **FLOATING
C1329 vin2.n64 vss 0.14fF $ **FLOATING
C1330 vin2.n65 vss 0.14fF $ **FLOATING
C1331 vin2.n66 vss 0.14fF $ **FLOATING
C1332 vin2.n67 vss 0.14fF $ **FLOATING
C1333 vin2.n68 vss 0.18fF $ **FLOATING
C1334 vin2.n69 vss 0.13fF $ **FLOATING
C1335 vin2.n70 vss 0.01fF $ **FLOATING
C1336 vin2.n71 vss 0.01fF $ **FLOATING
C1337 vin2.n72 vss 0.47fF $ **FLOATING
C1338 vin2.n73 vss 0.19fF $ **FLOATING
C1339 vin2.n74 vss 0.14fF $ **FLOATING
C1340 vin2.n75 vss 0.14fF $ **FLOATING
C1341 vin2.n76 vss 0.14fF $ **FLOATING
C1342 vin2.n77 vss 0.14fF $ **FLOATING
C1343 vin2.n78 vss 0.14fF $ **FLOATING
C1344 vin2.n79 vss 0.14fF $ **FLOATING
C1345 vin2.n80 vss 0.14fF $ **FLOATING
C1346 vin2.n81 vss 0.14fF $ **FLOATING
C1347 vin2.n82 vss 0.18fF $ **FLOATING
C1348 vin2.n83 vss 1.53fF $ **FLOATING
C1349 vin2.n84 vss 7.22fF $ **FLOATING
C1350 vout.n0 vss 0.07fF $ **FLOATING
C1351 vout.n1 vss 0.05fF $ **FLOATING
C1352 vout.t34 vss 6.87fF
C1353 vout.t33 vss 7.43fF
C1354 vout.t36 vss 6.11fF
C1355 vout.n2 vss 1.75fF $ **FLOATING
C1356 vout.t35 vss 9.40fF
C1357 vout.t0 vss 10.42fF
C1358 vout.t1 vss 5.74fF
C1359 vout.n3 vss 0.37fF $ **FLOATING
C1360 vout.n4 vss 0.37fF $ **FLOATING
C1361 vout.t3 vss 5.47fF
C1362 vout.n5 vss 1.52fF $ **FLOATING
C1363 vout.t2 vss 6.66fF
C1364 vout.n6 vss 3.10fF $ **FLOATING
C1365 pmos_3p3_CDNS_679510442370_0.S vss 3.68fF $ **FLOATING
C1366 vout.n7 vss 0.30fF $ **FLOATING
C1367 vout.n8 vss 0.17fF $ **FLOATING
C1368 vout.n9 vss 0.16fF $ **FLOATING
C1369 vout.n10 vss 0.30fF $ **FLOATING
C1370 vout.n11 vss 0.17fF $ **FLOATING
C1371 vout.n12 vss 5.60fF $ **FLOATING
C1372 vout.n13 vss 3.89fF $ **FLOATING
C1373 vout.n14 vss 3.24fF $ **FLOATING
C1374 vout.n15 vss 2.53fF $ **FLOATING
C1375 vout.n16 vss 0.01fF $ **FLOATING
C1376 vout.n17 vss 0.01fF $ **FLOATING
C1377 nmos_3p3_CDNS_679510442372_0.S vss 0.30fF $ **FLOATING
C1378 vout.n18 vss 0.05fF $ **FLOATING
C1379 vout.n19 vss 0.03fF $ **FLOATING
C1380 vout.n20 vss 0.03fF $ **FLOATING
C1381 vout.n21 vss 0.04fF $ **FLOATING
C1382 vout.n22 vss 0.04fF $ **FLOATING
C1383 vout.n23 vss 0.05fF $ **FLOATING
C1384 vout.n24 vss 0.01fF $ **FLOATING
C1385 vout.n25 vss 0.01fF $ **FLOATING
C1386 vout.n26 vss 0.01fF $ **FLOATING
C1387 vout.n27 vss 0.01fF $ **FLOATING
C1388 vout.n28 vss 0.56fF $ **FLOATING
C1389 vout.n29 vss 0.47fF $ **FLOATING
C1390 vout.n30 vss 0.05fF $ **FLOATING
C1391 vout.n31 vss 0.05fF $ **FLOATING
.ends


* File: opamp2_hspice.pex.netlist
* Created: Wed Mar 22 22:30:36 2023
* Program "Calibre xRC"
* Version "v2022.2_15.10"
* 
.include "opamp2_hspice.pex.netlist.pex"
.subckt opamp2_nodw  VBIASN VBIASP VDD VIN1 VIN2 VOUT VOUT_T VPROG VSS
* 
* VOUT_T	VOUT_T
* VBIASN	VBIASN
* VOUT	VOUT
* VBIASP	VBIASP
* VIN1	VIN1
* VIN2	VIN2
* VSS	VSS
* VPROG	VPROG
* VDD	VDD
XMMN25<4> N_VSS_MMN25<4>_d N_VSS_MMN25<4>_g N_VSS_MMN25<4>_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN25<3>@10 N_VSS_MMN25<3>@10_d N_VSS_MMN25<3>@10_g N_VSS_MMN25<3>@10_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN25<3>@9 N_VSS_MMN25<4>_s N_VSS_MMN25<3>@9_g N_VSS_MMN25<3>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@8 N_VSS_MMN25<3>@10_s N_VSS_MMN25<3>@8_g N_VSS_MMN25<3>@8_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@7 N_VSS_MMN25<3>@9_s N_VSS_MMN25<3>@7_g N_VSS_MMN25<3>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@6 N_VSS_MMN25<3>@8_s N_VSS_MMN25<3>@6_g N_VSS_MMN25<3>@6_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@5 N_VSS_MMN25<3>@7_s N_VSS_MMN25<3>@5_g N_VSS_MMN25<3>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@4 N_VSS_MMN25<3>@6_s N_VSS_MMN25<3>@4_g N_VSS_MMN25<3>@4_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@3 N_VSS_MMN25<3>@5_s N_VSS_MMN25<3>@3_g N_VSS_MMN25<3>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3>@2 N_VSS_MMN25<3>@4_s N_VSS_MMN25<3>@2_g N_VSS_MMN25<3>@2_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<3> N_VSS_MMN25<3>@3_s N_VSS_MMN25<3>_g N_VSS_MMN25<3>_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@10 N_VSS_MMN25<3>@2_s N_VSS_MMN25<2>@10_g N_VSS_MMN25<2>@10_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@9 N_VSS_MMN25<3>_s N_VSS_MMN25<2>@9_g N_VSS_MMN25<2>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@8 N_VSS_MMN25<2>@10_s N_VSS_MMN25<2>@8_g N_VSS_MMN25<2>@8_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@7 N_VSS_MMN25<2>@9_s N_VSS_MMN25<2>@7_g N_VSS_MMN25<2>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@6 N_VSS_MMN25<2>@8_s N_VSS_MMN25<2>@6_g N_VSS_MMN25<2>@6_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@5 N_VSS_MMN25<2>@7_s N_VSS_MMN25<2>@5_g N_VSS_MMN25<2>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@4 N_VSS_MMN25<2>@6_s N_VSS_MMN25<2>@4_g N_VSS_MMN25<2>@4_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@3 N_VSS_MMN25<2>@5_s N_VSS_MMN25<2>@3_g N_VSS_MMN25<2>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<2>@2 N_VSS_MMN25<2>@4_s N_VSS_MMN25<2>@2_g N_VSS_MMN25<2>@2_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN33 N_NET12_MMN33_d N_NET12_MMN33_g N_VSS_MMN33_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=4e-06 AD=1.04e-12 AS=1.76e-12 PD=4.52e-06 PS=8.88e-06 NRD=0.065
+ NRS=0.11 M=1 NF=1 PAR=1
XMMN34 N_VTAILN_MMN34_d N_NET12_MMN34_g N_VSS_MMN34_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=4e-06 AD=1.04e-12 AS=1.76e-12 PD=4.52e-06 PS=8.88e-06 NRD=0.065
+ NRS=0.11 M=1 NF=1 PAR=1
XMMN34@25 N_VTAILN_MMN34@25_d N_NET12_MMN34@25_g N_VSS_MMN34@25_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.76e-12 PD=4.52e-06
+ PS=8.88e-06 NRD=0.065 NRS=0.11 M=1 NF=1 PAR=1
XMMN30 N_NET8_MMN30_d N_NET8_MMN30_g N_NET12_MMN30_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2e-06 AD=8.8e-13 AS=5.2e-13 PD=4.88e-06 PS=2.52e-06 NRD=0.22
+ NRS=0.13 M=1 NF=1 PAR=1
XMMN30@10 N_NET8_MMN30@10_d N_NET8_MMN30@10_g N_NET12_MMN30@10_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=2e-06 AD=8.8e-13 AS=5.2e-13 PD=4.88e-06
+ PS=2.52e-06 NRD=0.22 NRS=0.13 M=1 NF=1 PAR=1
XMMN33@5 N_NET12_MMN33_d N_NET12_MMN33@5_g N_VSS_MMN33@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@24 N_VTAILN_MMN34_d N_NET12_MMN34@24_g N_VSS_MMN34@24_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@23 N_VTAILN_MMN34@25_d N_NET12_MMN34@23_g N_VSS_MMN34@23_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN30@9 N_NET8_MMN30@9_d N_NET8_MMN30@9_g N_NET12_MMN30_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN30@8 N_NET8_MMN30@8_d N_NET8_MMN30@8_g N_NET12_MMN30@10_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN33@4 N_NET12_MMN33@4_d N_NET12_MMN33@4_g N_VSS_MMN33@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@22 N_VTAILN_MMN34@22_d N_NET12_MMN34@22_g N_VSS_MMN34@24_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@21 N_VTAILN_MMN34@21_d N_NET12_MMN34@21_g N_VSS_MMN34@23_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN30@7 N_NET8_MMN30@9_d N_NET8_MMN30@7_g N_NET12_MMN30@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN30@6 N_NET8_MMN30@8_d N_NET8_MMN30@6_g N_NET12_MMN30@6_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN33@3 N_NET12_MMN33@4_d N_NET12_MMN33@3_g N_VSS_MMN33@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@20 N_VTAILN_MMN34@22_d N_NET12_MMN34@20_g N_VSS_MMN34@20_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@19 N_VTAILN_MMN34@21_d N_NET12_MMN34@19_g N_VSS_MMN34@19_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN30@5 N_NET8_MMN30@5_d N_NET8_MMN30@5_g N_NET12_MMN30@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN30@4 N_NET8_MMN30@4_d N_NET8_MMN30@4_g N_NET12_MMN30@6_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN33@2 N_NET12_MMN33@2_d N_NET12_MMN33@2_g N_VSS_MMN33@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.76e-12 AS=1.04e-12 PD=8.88e-06 PS=4.52e-06
+ NRD=0.11 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@18 N_VTAILN_MMN34@18_d N_NET12_MMN34@18_g N_VSS_MMN34@20_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.76e-12 AS=1.04e-12 PD=8.88e-06
+ PS=4.52e-06 NRD=0.11 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@17 N_VTAILN_MMN34@17_d N_NET12_MMN34@17_g N_VSS_MMN34@19_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.76e-12 AS=1.04e-12 PD=8.88e-06
+ PS=4.52e-06 NRD=0.11 NRS=0.065 M=1 NF=1 PAR=1
XMMN30@3 N_NET8_MMN30@5_d N_NET8_MMN30@3_g N_NET12_MMN30@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=8.8e-13 PD=2.52e-06 PS=4.88e-06
+ NRD=0.13 NRS=0.22 M=1 NF=1 PAR=1
XMMN30@2 N_NET8_MMN30@4_d N_NET8_MMN30@2_g N_NET12_MMN30@2_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=8.8e-13 PD=2.52e-06 PS=4.88e-06
+ NRD=0.13 NRS=0.22 M=1 NF=1 PAR=1
XMMN29 N_NET11_MMN29_d N_NET8_MMN29_g N_NET10_MMN29_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2.2e-07 AD=1.516e-13 AS=1.516e-13 PD=1.64e-06 PS=1.64e-06
+ NRD=3.13223 NRS=3.13223 M=1 NF=1 PAR=1
XMMN22 N_VSS_MMN22_d N_VSS_MMN22_g N_VSS_MMN22_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=4e-06 AD=1.76e-12 AS=1.76e-12 PD=8.88e-06 PS=8.88e-06 NRD=0.11
+ NRS=0.11 M=1 NF=1 PAR=1
XMMN32 N_NET9_MMN32_d N_NET9_MMN32_g N_VSS_MMN32_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN31 N_NET7_MMN31_d N_NET12_MMN31_g N_VSS_MMN31_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN35 N_NET10_MMN35_d N_NET12_MMN35_g N_VSS_MMN35_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN22@2 N_VSS_MMN22@2_d N_VSS_MMN22@2_g N_VSS_MMN22@2_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=5e-06 AD=2.2e-12 AS=2.2e-12 PD=1.088e-05 PS=1.088e-05
+ NRD=0.088 NRS=0.088 M=1 NF=1 PAR=1
XMMN34@16 N_VTAILN_MMN34@16_d N_NET12_MMN34@16_g N_VSS_MMN34@16_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.76e-12 PD=4.52e-06
+ PS=8.88e-06 NRD=0.065 NRS=0.11 M=1 NF=1 PAR=1
XMMN34@15 N_VTAILN_MMN34@15_d N_NET12_MMN34@15_g N_VSS_MMN34@15_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.76e-12 PD=4.52e-06
+ PS=8.88e-06 NRD=0.065 NRS=0.11 M=1 NF=1 PAR=1
XMMN34@14 N_VTAILN_MMN34@14_d N_NET12_MMN34@14_g N_VSS_MMN34@14_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.76e-12 PD=4.52e-06
+ PS=8.88e-06 NRD=0.065 NRS=0.11 M=1 NF=1 PAR=1
XMMN27 N_IABP_MMN27_d N_NET8_MMN27_g N_NET7_MMN27_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2e-06 AD=5.2e-13 AS=8.8e-13 PD=2.52e-06 PS=4.88e-06 NRD=0.13
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN28 N_IABN_MMN28_d N_IABN_MMN28_g N_NET9_MMN28_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=2e-06 AD=8.8e-13 AS=5.2e-13 PD=4.88e-06 PS=2.52e-06 NRD=0.22
+ NRS=0.13 M=1 NF=1 PAR=1
XMMN34@13 N_VTAILN_MMN34@16_d N_NET12_MMN34@13_g N_VSS_MMN34@13_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@12 N_VTAILN_MMN34@15_d N_NET12_MMN34@12_g N_VSS_MMN34@12_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@11 N_VTAILN_MMN34@14_d N_NET12_MMN34@11_g N_VSS_MMN34@11_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN27@5 N_IABP_MMN27_d N_NET8_MMN27@5_g N_NET7_MMN27@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN28@5 N_IABN_MMN28@5_d N_IABN_MMN28@5_g N_NET9_MMN28_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN34@10 N_VTAILN_MMN34@10_d N_NET12_MMN34@10_g N_VSS_MMN34@13_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06
+ PS=4.52e-06 NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@9 N_VTAILN_MMN34@9_d N_NET12_MMN34@9_g N_VSS_MMN34@12_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@8 N_VTAILN_MMN34@8_d N_NET12_MMN34@8_g N_VSS_MMN34@11_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN27@4 N_IABP_MMN27@4_d N_NET8_MMN27@4_g N_NET7_MMN27@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN28@4 N_IABN_MMN28@5_d N_IABN_MMN28@4_g N_NET9_MMN28@4_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN34@7 N_VTAILN_MMN34@10_d N_NET12_MMN34@7_g N_VSS_MMN34@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@6 N_VTAILN_MMN34@9_d N_NET12_MMN34@6_g N_VSS_MMN34@6_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@5 N_VTAILN_MMN34@8_d N_NET12_MMN34@5_g N_VSS_MMN34@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.04e-12 AS=1.04e-12 PD=4.52e-06 PS=4.52e-06
+ NRD=0.065 NRS=0.065 M=1 NF=1 PAR=1
XMMN27@3 N_IABP_MMN27@4_d N_NET8_MMN27@3_g N_NET7_MMN27@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN28@3 N_IABN_MMN28@3_d N_IABN_MMN28@3_g N_NET9_MMN28@4_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMN34@4 N_VTAILN_MMN34@4_d N_NET12_MMN34@4_g N_VSS_MMN34@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.76e-12 AS=1.04e-12 PD=8.88e-06 PS=4.52e-06
+ NRD=0.11 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@3 N_VTAILN_MMN34@3_d N_NET12_MMN34@3_g N_VSS_MMN34@6_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.76e-12 AS=1.04e-12 PD=8.88e-06 PS=4.52e-06
+ NRD=0.11 NRS=0.065 M=1 NF=1 PAR=1
XMMN34@2 N_VTAILN_MMN34@2_d N_NET12_MMN34@2_g N_VSS_MMN34@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=4e-06 AD=1.76e-12 AS=1.04e-12 PD=8.88e-06 PS=4.52e-06
+ NRD=0.11 NRS=0.065 M=1 NF=1 PAR=1
XMMN27@2 N_IABP_MMN27@2_d N_NET8_MMN27@2_g N_NET7_MMN27@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=8.8e-13 AS=5.2e-13 PD=4.88e-06 PS=2.52e-06
+ NRD=0.22 NRS=0.13 M=1 NF=1 PAR=1
XMMN28@2 N_IABN_MMN28@3_d N_IABN_MMN28@2_g N_NET9_MMN28@2_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=2e-06 AD=5.2e-13 AS=8.8e-13 PD=2.52e-06 PS=4.88e-06
+ NRD=0.13 NRS=0.22 M=1 NF=1 PAR=1
XMMN25<2> N_VSS_MMN25<2>_d N_VSS_MMN25<2>_g N_VSS_MMN25<2>_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN25<1>@10 N_VSS_MMN25<1>@10_d N_VSS_MMN25<1>@10_g N_VSS_MMN25<1>@10_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN25<1>@9 N_VSS_MMN25<2>_s N_VSS_MMN25<1>@9_g N_VSS_MMN25<1>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@8 N_VSS_MMN25<1>@10_s N_VSS_MMN25<1>@8_g N_VSS_MMN25<1>@8_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@7 N_VSS_MMN25<1>@9_s N_VSS_MMN25<1>@7_g N_VSS_MMN25<1>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@6 N_VSS_MMN25<1>@8_s N_VSS_MMN25<1>@6_g N_VSS_MMN25<1>@6_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@5 N_VSS_MMN25<1>@7_s N_VSS_MMN25<1>@5_g N_VSS_MMN25<1>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@4 N_VSS_MMN25<1>@6_s N_VSS_MMN25<1>@4_g N_VSS_MMN25<1>@4_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@3 N_VSS_MMN25<1>@5_s N_VSS_MMN25<1>@3_g N_VSS_MMN25<1>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1>@2 N_VSS_MMN25<1>@4_s N_VSS_MMN25<1>@2_g N_VSS_MMN25<1>@2_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<1> N_VSS_MMN25<1>@3_s N_VSS_MMN25<1>_g N_VSS_MMN25<1>_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@10 N_VSS_MMN25<1>@2_s N_VSS_MMN25<0>@10_g N_VSS_MMN25<0>@10_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@9 N_VSS_MMN25<1>_s N_VSS_MMN25<0>@9_g N_VSS_MMN25<0>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@8 N_VSS_MMN25<0>@10_s N_VSS_MMN25<0>@8_g N_VSS_MMN25<0>@8_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@7 N_VSS_MMN25<0>@9_s N_VSS_MMN25<0>@7_g N_VSS_MMN25<0>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@6 N_VSS_MMN25<0>@8_s N_VSS_MMN25<0>@6_g N_VSS_MMN25<0>@6_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@5 N_VSS_MMN25<0>@7_s N_VSS_MMN25<0>@5_g N_VSS_MMN25<0>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@4 N_VSS_MMN25<0>@6_s N_VSS_MMN25<0>@4_g N_VSS_MMN25<0>@4_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@3 N_VSS_MMN25<0>@5_s N_VSS_MMN25<0>@3_g N_VSS_MMN25<0>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0>@2 N_VSS_MMN25<0>@4_s N_VSS_MMN25<0>@2_g N_VSS_MMN25<0>@2_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3> N_NET4_MMN43<3>_d N_VIN2_MMN43<3>_g N_VTAILN_MMN43<3>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3> N_NET5_MMN42<3>_d N_VIN1_MMN42<3>_g N_VTAILN_MMN42<3>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@10 N_NET4_MMN43<2>@10_d N_VIN2_MMN43<2>@10_g N_VTAILN_MMN43<3>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@10 N_NET5_MMN42<2>@10_d N_VIN1_MMN42<2>@10_g N_VTAILN_MMN42<3>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@9 N_NET4_MMN43<2>@10_d N_VIN2_MMN43<2>@9_g N_VTAILN_MMN43<2>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@9 N_NET5_MMN42<2>@10_d N_VIN1_MMN42<2>@9_g N_VTAILN_MMN42<2>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@8 N_NET4_MMN43<2>@8_d N_VIN2_MMN43<2>@8_g N_VTAILN_MMN43<2>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@8 N_NET5_MMN42<2>@8_d N_VIN1_MMN42<2>@8_g N_VTAILN_MMN42<2>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@7 N_NET4_MMN43<2>@8_d N_VIN2_MMN43<2>@7_g N_VTAILN_MMN43<2>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@7 N_NET5_MMN42<2>@8_d N_VIN1_MMN42<2>@7_g N_VTAILN_MMN42<2>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@6 N_NET4_MMN43<2>@6_d N_VIN2_MMN43<2>@6_g N_VTAILN_MMN43<2>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@6 N_NET5_MMN42<2>@6_d N_VIN1_MMN42<2>@6_g N_VTAILN_MMN42<2>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@5 N_NET4_MMN43<2>@6_d N_VIN2_MMN43<2>@5_g N_VTAILN_MMN43<2>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@5 N_NET5_MMN42<2>@6_d N_VIN1_MMN42<2>@5_g N_VTAILN_MMN42<2>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@4 N_NET4_MMN43<2>@4_d N_VIN2_MMN43<2>@4_g N_VTAILN_MMN43<2>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@4 N_NET5_MMN42<2>@4_d N_VIN1_MMN42<2>@4_g N_VTAILN_MMN42<2>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@3 N_NET4_MMN43<2>@4_d N_VIN2_MMN43<2>@3_g N_VTAILN_MMN43<2>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@3 N_NET5_MMN42<2>@4_d N_VIN1_MMN42<2>@3_g N_VTAILN_MMN42<2>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2>@2 N_NET4_MMN43<2>@2_d N_VIN2_MMN43<2>@2_g N_VTAILN_MMN43<2>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2>@2 N_NET5_MMN42<2>@2_d N_VIN1_MMN42<2>@2_g N_VTAILN_MMN42<2>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<2> N_NET5_MMN42<2>_d N_VIN1_MMN42<2>_g N_VTAILN_MMN42<2>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<2> N_NET4_MMN43<2>_d N_VIN2_MMN43<2>_g N_VTAILN_MMN43<2>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@10 N_NET5_MMN42<1>@10_d N_VIN1_MMN42<1>@10_g N_VTAILN_MMN42<2>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@10 N_NET4_MMN43<1>@10_d N_VIN2_MMN43<1>@10_g N_VTAILN_MMN43<2>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@9 N_NET5_MMN42<1>@10_d N_VIN1_MMN42<1>@9_g N_VTAILN_MMN42<1>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@9 N_NET4_MMN43<1>@10_d N_VIN2_MMN43<1>@9_g N_VTAILN_MMN43<1>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@8 N_NET5_MMN42<1>@8_d N_VIN1_MMN42<1>@8_g N_VTAILN_MMN42<1>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@8 N_NET4_MMN43<1>@8_d N_VIN2_MMN43<1>@8_g N_VTAILN_MMN43<1>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@7 N_NET5_MMN42<1>@8_d N_VIN1_MMN42<1>@7_g N_VTAILN_MMN42<1>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@7 N_NET4_MMN43<1>@8_d N_VIN2_MMN43<1>@7_g N_VTAILN_MMN43<1>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@6 N_NET5_MMN42<1>@6_d N_VIN1_MMN42<1>@6_g N_VTAILN_MMN42<1>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@6 N_NET4_MMN43<1>@6_d N_VIN2_MMN43<1>@6_g N_VTAILN_MMN43<1>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@5 N_NET5_MMN42<1>@6_d N_VIN1_MMN42<1>@5_g N_VTAILN_MMN42<1>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@5 N_NET4_MMN43<1>@6_d N_VIN2_MMN43<1>@5_g N_VTAILN_MMN43<1>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@4 N_NET5_MMN42<1>@4_d N_VIN1_MMN42<1>@4_g N_VTAILN_MMN42<1>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@4 N_NET4_MMN43<1>@4_d N_VIN2_MMN43<1>@4_g N_VTAILN_MMN43<1>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@3 N_NET5_MMN42<1>@4_d N_VIN1_MMN42<1>@3_g N_VTAILN_MMN42<1>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@3 N_NET4_MMN43<1>@4_d N_VIN2_MMN43<1>@3_g N_VTAILN_MMN43<1>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1>@2 N_NET5_MMN42<1>@2_d N_VIN1_MMN42<1>@2_g N_VTAILN_MMN42<1>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1>@2 N_NET4_MMN43<1>@2_d N_VIN2_MMN43<1>@2_g N_VTAILN_MMN43<1>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<1> N_NET5_MMN42<1>_d N_VIN1_MMN42<1>_g N_VTAILN_MMN42<1>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<1> N_NET4_MMN43<1>_d N_VIN2_MMN43<1>_g N_VTAILN_MMN43<1>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@10 N_NET5_MMN42<0>@10_d N_VIN1_MMN42<0>@10_g N_VTAILN_MMN42<1>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@10 N_NET4_MMN43<0>@10_d N_VIN2_MMN43<0>@10_g N_VTAILN_MMN43<1>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@9 N_NET5_MMN42<0>@10_d N_VIN1_MMN42<0>@9_g N_VTAILN_MMN42<0>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@9 N_NET4_MMN43<0>@10_d N_VIN2_MMN43<0>@9_g N_VTAILN_MMN43<0>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@8 N_NET5_MMN42<0>@8_d N_VIN1_MMN42<0>@8_g N_VTAILN_MMN42<0>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@8 N_NET4_MMN43<0>@8_d N_VIN2_MMN43<0>@8_g N_VTAILN_MMN43<0>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@7 N_NET5_MMN42<0>@8_d N_VIN1_MMN42<0>@7_g N_VTAILN_MMN42<0>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@7 N_NET4_MMN43<0>@8_d N_VIN2_MMN43<0>@7_g N_VTAILN_MMN43<0>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@6 N_NET5_MMN42<0>@6_d N_VIN1_MMN42<0>@6_g N_VTAILN_MMN42<0>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@6 N_NET4_MMN43<0>@6_d N_VIN2_MMN43<0>@6_g N_VTAILN_MMN43<0>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@5 N_NET5_MMN42<0>@6_d N_VIN1_MMN42<0>@5_g N_VTAILN_MMN42<0>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@5 N_NET4_MMN43<0>@6_d N_VIN2_MMN43<0>@5_g N_VTAILN_MMN43<0>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@4 N_NET5_MMN42<0>@4_d N_VIN1_MMN42<0>@4_g N_VTAILN_MMN42<0>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@4 N_NET4_MMN43<0>@4_d N_VIN2_MMN43<0>@4_g N_VTAILN_MMN43<0>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@3 N_NET5_MMN42<0>@4_d N_VIN1_MMN42<0>@3_g N_VTAILN_MMN42<0>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@3 N_NET4_MMN43<0>@4_d N_VIN2_MMN43<0>@3_g N_VTAILN_MMN43<0>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0>@2 N_NET5_MMN42<0>@2_d N_VIN1_MMN42<0>@2_g N_VTAILN_MMN42<0>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0>@2 N_NET4_MMN43<0>@2_d N_VIN2_MMN43<0>@2_g N_VTAILN_MMN43<0>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<0> N_NET4_MMN43<0>_d N_VIN2_MMN43<0>_g N_VTAILN_MMN43<0>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<0> N_NET5_MMN42<0>_d N_VIN1_MMN42<0>_g N_VTAILN_MMN42<0>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@10 N_NET4_MMN43<3>@10_d N_VIN2_MMN43<3>@10_g N_VTAILN_MMN43<0>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@10 N_NET5_MMN42<3>@10_d N_VIN1_MMN42<3>@10_g N_VTAILN_MMN42<0>_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@9 N_NET4_MMN43<3>@10_d N_VIN2_MMN43<3>@9_g N_VTAILN_MMN43<3>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@9 N_NET5_MMN42<3>@10_d N_VIN1_MMN42<3>@9_g N_VTAILN_MMN42<3>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@8 N_NET4_MMN43<3>@8_d N_VIN2_MMN43<3>@8_g N_VTAILN_MMN43<3>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@8 N_NET5_MMN42<3>@8_d N_VIN1_MMN42<3>@8_g N_VTAILN_MMN42<3>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@7 N_NET4_MMN43<3>@8_d N_VIN2_MMN43<3>@7_g N_VTAILN_MMN43<3>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@7 N_NET5_MMN42<3>@8_d N_VIN1_MMN42<3>@7_g N_VTAILN_MMN42<3>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@6 N_NET4_MMN43<3>@6_d N_VIN2_MMN43<3>@6_g N_VTAILN_MMN43<3>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@6 N_NET5_MMN42<3>@6_d N_VIN1_MMN42<3>@6_g N_VTAILN_MMN42<3>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@5 N_NET4_MMN43<3>@6_d N_VIN2_MMN43<3>@5_g N_VTAILN_MMN43<3>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@5 N_NET5_MMN42<3>@6_d N_VIN1_MMN42<3>@5_g N_VTAILN_MMN42<3>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@4 N_NET4_MMN43<3>@4_d N_VIN2_MMN43<3>@4_g N_VTAILN_MMN43<3>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@4 N_NET5_MMN42<3>@4_d N_VIN1_MMN42<3>@4_g N_VTAILN_MMN42<3>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@3 N_NET4_MMN43<3>@4_d N_VIN2_MMN43<3>@3_g N_VTAILN_MMN43<3>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@3 N_NET5_MMN42<3>@4_d N_VIN1_MMN42<3>@3_g N_VTAILN_MMN42<3>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN43<3>@2 N_NET4_MMN43<3>@2_d N_VIN2_MMN43<3>@2_g N_VTAILN_MMN43<3>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN42<3>@2 N_NET5_MMN42<3>@2_d N_VIN1_MMN42<3>@2_g N_VTAILN_MMN42<3>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<0> N_VSS_MMN25<0>_d N_VSS_MMN25<0>_g N_VSS_MMN25<0>_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN40 N_VOUT_MMN40_d N_NET6_MMN40_g N_VSS_MMN40_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05 NRD=0.044
+ NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@10 N_VSS_MMN25<0>_s N_VSS_MMN25<4>@10_g N_VSS_MMN25<4>@10_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@10 N_VOUT_MMN40@10_d N_NET6_MMN40@10_g N_VSS_MMN40_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@9 N_VSS_MMN25<4>@10_s N_VSS_MMN25<4>@9_g N_VSS_MMN25<4>@9_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@9 N_VOUT_MMN40@10_d N_NET6_MMN40@9_g N_VSS_MMN40@9_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@8 N_VSS_MMN25<4>@9_s N_VSS_MMN25<4>@8_g N_VSS_MMN25<4>@8_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@8 N_VOUT_MMN40@8_d N_NET6_MMN40@8_g N_VSS_MMN40@9_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@7 N_VSS_MMN25<4>@8_s N_VSS_MMN25<4>@7_g N_VSS_MMN25<4>@7_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@7 N_VOUT_MMN40@8_d N_NET6_MMN40@7_g N_VSS_MMN40@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@6 N_VSS_MMN25<4>@7_s N_VSS_MMN25<4>@6_g N_VSS_MMN25<4>@6_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@6 N_VOUT_MMN40@6_d N_NET6_MMN40@6_g N_VSS_MMN40@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@5 N_VSS_MMN25<4>@6_s N_VSS_MMN25<4>@5_g N_VSS_MMN25<4>@5_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@5 N_VOUT_MMN40@6_d N_NET6_MMN40@5_g N_VSS_MMN40@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@4 N_VSS_MMN25<4>@5_s N_VSS_MMN25<4>@4_g N_VSS_MMN25<4>@4_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@4 N_VOUT_MMN40@4_d N_NET6_MMN40@4_g N_VSS_MMN40@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@3 N_VSS_MMN25<4>@4_s N_VSS_MMN25<4>@3_g N_VSS_MMN25<4>@3_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@3 N_VOUT_MMN40@4_d N_NET6_MMN40@3_g N_VSS_MMN40@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN25<4>@2 N_VSS_MMN25<4>@3_s N_VSS_MMN25<4>@2_g N_VSS_MMN25<4>@2_s
+ N_VSS_MMN25<4>_b NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN40@2 N_VOUT_MMN40@2_d N_NET6_MMN40@2_g N_VSS_MMN40@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05
+ NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN44 N_NET1_MMN44_d N_IABN_MMN44_g N_NET6_MMN44_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=1e-05 AD=4.4e-12 AS=4.4e-12 PD=2.088e-05 PS=2.088e-05 NRD=0.044
+ NRS=0.044 M=1 NF=1 PAR=1
XMMN41 N_NET3_MMN41_d N_IABN_MMN41_g N_NET2_MMN41_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=1e-05 AD=4.4e-12 AS=4.4e-12 PD=2.088e-05 PS=2.088e-05 NRD=0.044
+ NRS=0.044 M=1 NF=1 PAR=1
XMMN36 N_NET13_MMN36_d N_NET2_MMN36_g N_VSS_MMN36_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05 NRD=0.026
+ NRS=0.044 M=1 NF=1 PAR=1
XMMN38 N_NET2_MMN38_d N_VBIASN_MMN38_g N_NET13_MMN38_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05 NRD=0.044
+ NRS=0.026 M=1 NF=1 PAR=1
XMMN36@2 N_NET13_MMN36_d N_NET2_MMN36@2_g N_VSS_MMN36@2_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN38@2 N_NET2_MMN38@2_d N_VBIASN_MMN38@2_g N_NET13_MMN38_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05
+ NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN37 N_NET14_MMN37_d N_NET2_MMN37_g N_VSS_MMN37_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05 NRD=0.026
+ NRS=0.044 M=1 NF=1 PAR=1
XMMN39 N_NET6_MMN39_d N_VBIASN_MMN39_g N_NET14_MMN39_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=1e-06 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05 NRD=0.044
+ NRS=0.026 M=1 NF=1 PAR=1
XMMN37@2 N_NET14_MMN37_d N_NET2_MMN37@2_g N_VSS_MMN37@2_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN39@2 N_NET6_MMN39@2_d N_VBIASN_MMN39@2_g N_NET14_MMN39_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=1e-06 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05
+ NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN3 N_VOUT_T_MMN3_d N_VDD_MMN3_g N_VOUT_MMN3_s N_VSS_MMN25<4>_b NMOS_3P3
+ L=2.8e-07 W=1e-06 AD=4.4e-13 AS=2.6e-13 PD=2.88e-06 PS=1.52e-06 NRD=0.44
+ NRS=0.26 M=1 NF=1 PAR=1
XMMN3@12 N_VOUT_T_MMN3@12_d N_VDD_MMN3@12_g N_VOUT_MMN3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@11 N_VOUT_T_MMN3@12_d N_VDD_MMN3@11_g N_VOUT_MMN3@11_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@10 N_VOUT_T_MMN3@10_d N_VDD_MMN3@10_g N_VOUT_MMN3@11_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@9 N_VOUT_T_MMN3@10_d N_VDD_MMN3@9_g N_VOUT_MMN3@9_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@8 N_VOUT_T_MMN3@8_d N_VDD_MMN3@8_g N_VOUT_MMN3@9_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@7 N_VOUT_T_MMN3@8_d N_VDD_MMN3@7_g N_VOUT_MMN3@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@6 N_VOUT_T_MMN3@6_d N_VDD_MMN3@6_g N_VOUT_MMN3@7_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@5 N_VOUT_T_MMN3@6_d N_VDD_MMN3@5_g N_VOUT_MMN3@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@4 N_VOUT_T_MMN3@4_d N_VDD_MMN3@4_g N_VOUT_MMN3@5_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@3 N_VOUT_T_MMN3@4_d N_VDD_MMN3@3_g N_VOUT_MMN3@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=2.6e-13 AS=2.6e-13 PD=1.52e-06 PS=1.52e-06
+ NRD=0.26 NRS=0.26 M=1 NF=1 PAR=1
XMMN3@2 N_VOUT_T_MMN3@2_d N_VDD_MMN3@2_g N_VOUT_MMN3@3_s N_VSS_MMN25<4>_b
+ NMOS_3P3 L=2.8e-07 W=1e-06 AD=4.4e-13 AS=2.6e-13 PD=2.88e-06 PS=1.52e-06
+ NRD=0.44 NRS=0.26 M=1 NF=1 PAR=1
XMMN23 N_VDD_MMN23_d N_VDD_MMN23_g N_VDD_MMN23_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN23@18 N_VDD_MMN23@18_d N_VDD_MMN23@18_g N_VDD_MMN23@18_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06
+ NRD=0.22 NRS=0.22 M=1 NF=1 PAR=1
XMMN24 N_VDD_MMN24_d N_VDD_MMN24_g N_VDD_MMN24_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06 NRD=0.176
+ NRS=0.176 M=1 NF=1 PAR=1
XMMN24@18 N_VDD_MMN24@18_d N_VDD_MMN24@18_g N_VDD_MMN24@18_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@17 N_VDD_MMN24@17_d N_VDD_MMN24@17_g N_VDD_MMN24@17_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@16 N_VDD_MMN24@16_d N_VDD_MMN24@16_g N_VDD_MMN24@16_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@15 N_VDD_MMN24@15_d N_VDD_MMN24@15_g N_VDD_MMN24@15_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@14 N_VDD_MMN24@14_d N_VDD_MMN24@14_g N_VDD_MMN24@14_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@13 N_VDD_MMN24@13_d N_VDD_MMN24@13_g N_VDD_MMN24@13_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP25 N_IABP_MMP25_d N_IABP_MMP25_g N_NET17_MMP25_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06 NRD=0.176
+ NRS=0.176 M=1 NF=1 PAR=1
XMMP25@4 N_IABP_MMP25@4_d N_IABP_MMP25@4_g N_NET17_MMP25@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@12 N_VDD_MMN24@12_d N_VDD_MMN24@12_g N_VDD_MMN24@12_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@11 N_VDD_MMN24@11_d N_VDD_MMN24@11_g N_VDD_MMN24@11_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@10 N_VDD_MMN24@10_d N_VDD_MMN24@10_g N_VDD_MMN24@10_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP30 N_NET17_MMP30_d N_NET17_MMP30_g N_VDD_MMP30_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMP26 N_NET8_MMP26_d N_VPROG_MMP26_g N_VDD_MMP26_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN24@9 N_VDD_MMN24@9_d N_VDD_MMN24@9_g N_VDD_MMN24@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP25@3 N_IABP_MMP25@3_d N_IABP_MMP25@3_g N_NET17_MMP25@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP25@2 N_IABP_MMP25@2_d N_IABP_MMP25@2_g N_NET17_MMP25@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@8 N_VDD_MMN24@8_d N_VDD_MMN24@8_g N_VDD_MMN24@8_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@7 N_VDD_MMN24@7_d N_VDD_MMN24@7_g N_VDD_MMN24@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@6 N_VDD_MMN24@6_d N_VDD_MMN24@6_g N_VDD_MMN24@6_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@5 N_VDD_MMN24@5_d N_VDD_MMN24@5_g N_VDD_MMN24@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP24 N_IABN_MMP24_d N_NET11_MMP24_g N_NET16_MMP24_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06 NRD=0.176
+ NRS=0.176 M=1 NF=1 PAR=1
XMMP24@4 N_IABN_MMP24@4_d N_NET11_MMP24@4_g N_NET16_MMP24@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP23 N_NET11_MMP23_d N_NET11_MMP23_g N_NET15_MMP23_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06 NRD=0.176
+ NRS=0.176 M=1 NF=1 PAR=1
XMMP23@4 N_NET11_MMP23@4_d N_NET11_MMP23@4_g N_NET15_MMP23@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@4 N_VDD_MMN24@4_d N_VDD_MMN24@4_g N_VDD_MMN24@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP29 N_NET16_MMP29_d N_NET15_MMP29_g N_VDD_MMP29_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMP28 N_NET15_MMP28_d N_NET15_MMP28_g N_VDD_MMP28_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=2e-06 AD=8.8e-13 AS=8.8e-13 PD=4.88e-06 PS=4.88e-06 NRD=0.22
+ NRS=0.22 M=1 NF=1 PAR=1
XMMN24@3 N_VDD_MMN24@3_d N_VDD_MMN24@3_g N_VDD_MMN24@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP24@3 N_IABN_MMP24@3_d N_NET11_MMP24@3_g N_NET16_MMP24@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP24@2 N_IABN_MMP24@2_d N_NET11_MMP24@2_g N_NET16_MMP24@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP23@3 N_NET11_MMP23@3_d N_NET11_MMP23@3_g N_NET15_MMP23@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP23@2 N_NET11_MMP23@2_d N_NET11_MMP23@2_g N_NET15_MMP23@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN24@2 N_VDD_MMN24@2_d N_VDD_MMN24@2_g N_VDD_MMN24@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=1e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@17 N_VDD_MMN23@17_d N_VDD_MMN23@17_g N_VDD_MMN23@17_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27 N_VTAILP_MMP27_d N_NET15_MMP27_g N_VDD_MMP27_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06 NRD=0.176
+ NRS=0.176 M=1 NF=1 PAR=1
XMMP27@40 N_VTAILP_MMP27@40_d N_NET15_MMP27@40_g N_VDD_MMP27@40_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@39 N_VTAILP_MMP27@39_d N_NET15_MMP27@39_g N_VDD_MMP27@39_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@38 N_VTAILP_MMP27@38_d N_NET15_MMP27@38_g N_VDD_MMP27@38_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@37 N_VTAILP_MMP27@37_d N_NET15_MMP27@37_g N_VDD_MMP27@37_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@36 N_VTAILP_MMP27@36_d N_NET15_MMP27@36_g N_VDD_MMP27@36_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@16 N_VDD_MMN23@16_d N_VDD_MMN23@16_g N_VDD_MMN23@16_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@15 N_VDD_MMN23@15_d N_VDD_MMN23@15_g N_VDD_MMN23@15_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@35 N_VTAILP_MMP27@35_d N_NET15_MMP27@35_g N_VDD_MMP27@35_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@34 N_VTAILP_MMP27@34_d N_NET15_MMP27@34_g N_VDD_MMP27@34_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@33 N_VTAILP_MMP27@33_d N_NET15_MMP27@33_g N_VDD_MMP27@33_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@32 N_VTAILP_MMP27@32_d N_NET15_MMP27@32_g N_VDD_MMP27@32_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@31 N_VTAILP_MMP27@31_d N_NET15_MMP27@31_g N_VDD_MMP27@31_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@30 N_VTAILP_MMP27@30_d N_NET15_MMP27@30_g N_VDD_MMP27@30_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@14 N_VDD_MMN23@14_d N_VDD_MMN23@14_g N_VDD_MMN23@14_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@13 N_VDD_MMN23@13_d N_VDD_MMN23@13_g N_VDD_MMN23@13_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@29 N_VTAILP_MMP27@29_d N_NET15_MMP27@29_g N_VDD_MMP27@29_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@28 N_VTAILP_MMP27@28_d N_NET15_MMP27@28_g N_VDD_MMP27@28_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@27 N_VTAILP_MMP27@27_d N_NET15_MMP27@27_g N_VDD_MMP27@27_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@26 N_VTAILP_MMP27@26_d N_NET15_MMP27@26_g N_VDD_MMP27@26_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@25 N_VTAILP_MMP27@25_d N_NET15_MMP27@25_g N_VDD_MMP27@25_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@24 N_VTAILP_MMP27@24_d N_NET15_MMP27@24_g N_VDD_MMP27@24_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@12 N_VDD_MMN23@12_d N_VDD_MMN23@12_g N_VDD_MMN23@12_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@11 N_VDD_MMN23@11_d N_VDD_MMN23@11_g N_VDD_MMN23@11_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@23 N_VTAILP_MMP27@23_d N_NET15_MMP27@23_g N_VDD_MMP27@23_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@22 N_VTAILP_MMP27@22_d N_NET15_MMP27@22_g N_VDD_MMP27@22_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@21 N_VTAILP_MMP27@21_d N_NET15_MMP27@21_g N_VDD_MMP27@21_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@20 N_VTAILP_MMP27@20_d N_NET15_MMP27@20_g N_VDD_MMP27@20_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@19 N_VTAILP_MMP27@19_d N_NET15_MMP27@19_g N_VDD_MMP27@19_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@18 N_VTAILP_MMP27@18_d N_NET15_MMP27@18_g N_VDD_MMP27@18_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@10 N_VDD_MMN23@10_d N_VDD_MMN23@10_g N_VDD_MMN23@10_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@9 N_VDD_MMN23@9_d N_VDD_MMN23@9_g N_VDD_MMN23@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@17 N_VTAILP_MMP27@17_d N_NET15_MMP27@17_g N_VDD_MMP27@17_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@16 N_VTAILP_MMP27@16_d N_NET15_MMP27@16_g N_VDD_MMP27@16_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@15 N_VTAILP_MMP27@15_d N_NET15_MMP27@15_g N_VDD_MMP27@15_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@14 N_VTAILP_MMP27@14_d N_NET15_MMP27@14_g N_VDD_MMP27@14_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@13 N_VTAILP_MMP27@13_d N_NET15_MMP27@13_g N_VDD_MMP27@13_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@12 N_VTAILP_MMP27@12_d N_NET15_MMP27@12_g N_VDD_MMP27@12_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@8 N_VDD_MMN23@8_d N_VDD_MMN23@8_g N_VDD_MMN23@8_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@7 N_VDD_MMN23@7_d N_VDD_MMN23@7_g N_VDD_MMN23@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@11 N_VTAILP_MMP27@11_d N_NET15_MMP27@11_g N_VDD_MMP27@11_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@10 N_VTAILP_MMP27@10_d N_NET15_MMP27@10_g N_VDD_MMP27@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06
+ PS=5.88e-06 NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@9 N_VTAILP_MMP27@9_d N_NET15_MMP27@9_g N_VDD_MMP27@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@8 N_VTAILP_MMP27@8_d N_NET15_MMP27@8_g N_VDD_MMP27@8_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@7 N_VTAILP_MMP27@7_d N_NET15_MMP27@7_g N_VDD_MMP27@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@6 N_VTAILP_MMP27@6_d N_NET15_MMP27@6_g N_VDD_MMP27@6_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@6 N_VDD_MMN23@6_d N_VDD_MMN23@6_g N_VDD_MMN23@6_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@5 N_VDD_MMN23@5_d N_VDD_MMN23@5_g N_VDD_MMN23@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@4 N_VDD_MMN23@4_d N_VDD_MMN23@4_g N_VDD_MMN23@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@5 N_VTAILP_MMP27@5_d N_NET15_MMP27@5_g N_VDD_MMP27@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@4 N_VTAILP_MMP27@4_d N_NET15_MMP27@4_g N_VDD_MMP27@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@3 N_VTAILP_MMP27@3_d N_NET15_MMP27@3_g N_VDD_MMP27@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP27@2 N_VTAILP_MMP27@2_d N_NET15_MMP27@2_g N_VDD_MMP27@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@3 N_VDD_MMN23@3_d N_VDD_MMN23@3_g N_VDD_MMN23@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMN23@2 N_VDD_MMN23@2_d N_VDD_MMN23@2_g N_VDD_MMN23@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=2.5e-06 AD=1.1e-12 AS=1.1e-12 PD=5.88e-06 PS=5.88e-06
+ NRD=0.176 NRS=0.176 M=1 NF=1 PAR=1
XMMP22<3> N_NET14_MMP22<3>_d N_VIN2_MMP22<3>_g N_VTAILP_MMP22<3>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<3> N_NET13_MMP21<3>_d N_VIN1_MMP21<3>_g N_VTAILP_MMP21<3>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<2>@10 N_NET14_MMP22<3>_d N_VIN2_MMP22<2>@10_g N_VTAILP_MMP22<2>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@10 N_NET13_MMP21<3>_d N_VIN1_MMP21<2>@10_g N_VTAILP_MMP21<2>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@9 N_NET14_MMP22<2>@9_d N_VIN2_MMP22<2>@9_g N_VTAILP_MMP22<2>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@9 N_NET13_MMP21<2>@9_d N_VIN1_MMP21<2>@9_g N_VTAILP_MMP21<2>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@8 N_NET14_MMP22<2>@9_d N_VIN2_MMP22<2>@8_g N_VTAILP_MMP22<2>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@8 N_NET13_MMP21<2>@9_d N_VIN1_MMP21<2>@8_g N_VTAILP_MMP21<2>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@7 N_NET14_MMP22<2>@7_d N_VIN2_MMP22<2>@7_g N_VTAILP_MMP22<2>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@7 N_NET13_MMP21<2>@7_d N_VIN1_MMP21<2>@7_g N_VTAILP_MMP21<2>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@6 N_NET14_MMP22<2>@7_d N_VIN2_MMP22<2>@6_g N_VTAILP_MMP22<2>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@6 N_NET13_MMP21<2>@7_d N_VIN1_MMP21<2>@6_g N_VTAILP_MMP21<2>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@5 N_NET14_MMP22<2>@5_d N_VIN2_MMP22<2>@5_g N_VTAILP_MMP22<2>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@5 N_NET13_MMP21<2>@5_d N_VIN1_MMP21<2>@5_g N_VTAILP_MMP21<2>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@4 N_NET14_MMP22<2>@5_d N_VIN2_MMP22<2>@4_g N_VTAILP_MMP22<2>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@4 N_NET13_MMP21<2>@5_d N_VIN1_MMP21<2>@4_g N_VTAILP_MMP21<2>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@3 N_NET14_MMP22<2>@3_d N_VIN2_MMP22<2>@3_g N_VTAILP_MMP22<2>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<2>@3 N_NET13_MMP21<2>@3_d N_VIN1_MMP21<2>@3_g N_VTAILP_MMP21<2>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<2>@2 N_NET14_MMP22<2>@3_d N_VIN2_MMP22<2>@2_g N_VTAILP_MMP22<2>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<2>@2 N_NET13_MMP21<2>@3_d N_VIN1_MMP21<2>@2_g N_VTAILP_MMP21<2>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<2> N_NET13_MMP21<2>_d N_VIN1_MMP21<2>_g N_VTAILP_MMP21<2>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<2> N_NET14_MMP22<2>_d N_VIN2_MMP22<2>_g N_VTAILP_MMP22<2>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<1>@10 N_NET13_MMP21<2>_d N_VIN1_MMP21<1>@10_g N_VTAILP_MMP21<1>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@10 N_NET14_MMP22<2>_d N_VIN2_MMP22<1>@10_g N_VTAILP_MMP22<1>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@9 N_NET13_MMP21<1>@9_d N_VIN1_MMP21<1>@9_g N_VTAILP_MMP21<1>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@9 N_NET14_MMP22<1>@9_d N_VIN2_MMP22<1>@9_g N_VTAILP_MMP22<1>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@8 N_NET13_MMP21<1>@9_d N_VIN1_MMP21<1>@8_g N_VTAILP_MMP21<1>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@8 N_NET14_MMP22<1>@9_d N_VIN2_MMP22<1>@8_g N_VTAILP_MMP22<1>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@7 N_NET13_MMP21<1>@7_d N_VIN1_MMP21<1>@7_g N_VTAILP_MMP21<1>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@7 N_NET14_MMP22<1>@7_d N_VIN2_MMP22<1>@7_g N_VTAILP_MMP22<1>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@6 N_NET13_MMP21<1>@7_d N_VIN1_MMP21<1>@6_g N_VTAILP_MMP21<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@6 N_NET14_MMP22<1>@7_d N_VIN2_MMP22<1>@6_g N_VTAILP_MMP22<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@5 N_NET13_MMP21<1>@5_d N_VIN1_MMP21<1>@5_g N_VTAILP_MMP21<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@5 N_NET14_MMP22<1>@5_d N_VIN2_MMP22<1>@5_g N_VTAILP_MMP22<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@4 N_NET13_MMP21<1>@5_d N_VIN1_MMP21<1>@4_g N_VTAILP_MMP21<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@4 N_NET14_MMP22<1>@5_d N_VIN2_MMP22<1>@4_g N_VTAILP_MMP22<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@3 N_NET13_MMP21<1>@3_d N_VIN1_MMP21<1>@3_g N_VTAILP_MMP21<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<1>@3 N_NET14_MMP22<1>@3_d N_VIN2_MMP22<1>@3_g N_VTAILP_MMP22<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<1>@2 N_NET13_MMP21<1>@3_d N_VIN1_MMP21<1>@2_g N_VTAILP_MMP21<1>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<1>@2 N_NET14_MMP22<1>@3_d N_VIN2_MMP22<1>@2_g N_VTAILP_MMP22<1>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<1> N_NET13_MMP21<1>_d N_VIN1_MMP21<1>_g N_VTAILP_MMP21<1>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<1> N_NET14_MMP22<1>_d N_VIN2_MMP22<1>_g N_VTAILP_MMP22<1>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<0>@10 N_NET13_MMP21<1>_d N_VIN1_MMP21<0>@10_g N_VTAILP_MMP21<0>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@10 N_NET14_MMP22<1>_d N_VIN2_MMP22<0>@10_g N_VTAILP_MMP22<0>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@9 N_NET13_MMP21<0>@9_d N_VIN1_MMP21<0>@9_g N_VTAILP_MMP21<0>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@9 N_NET14_MMP22<0>@9_d N_VIN2_MMP22<0>@9_g N_VTAILP_MMP22<0>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@8 N_NET13_MMP21<0>@9_d N_VIN1_MMP21<0>@8_g N_VTAILP_MMP21<0>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@8 N_NET14_MMP22<0>@9_d N_VIN2_MMP22<0>@8_g N_VTAILP_MMP22<0>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@7 N_NET13_MMP21<0>@7_d N_VIN1_MMP21<0>@7_g N_VTAILP_MMP21<0>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@7 N_NET14_MMP22<0>@7_d N_VIN2_MMP22<0>@7_g N_VTAILP_MMP22<0>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@6 N_NET13_MMP21<0>@7_d N_VIN1_MMP21<0>@6_g N_VTAILP_MMP21<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@6 N_NET14_MMP22<0>@7_d N_VIN2_MMP22<0>@6_g N_VTAILP_MMP22<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@5 N_NET13_MMP21<0>@5_d N_VIN1_MMP21<0>@5_g N_VTAILP_MMP21<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@5 N_NET14_MMP22<0>@5_d N_VIN2_MMP22<0>@5_g N_VTAILP_MMP22<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@4 N_NET13_MMP21<0>@5_d N_VIN1_MMP21<0>@4_g N_VTAILP_MMP21<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@4 N_NET14_MMP22<0>@5_d N_VIN2_MMP22<0>@4_g N_VTAILP_MMP22<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@3 N_NET13_MMP21<0>@3_d N_VIN1_MMP21<0>@3_g N_VTAILP_MMP21<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<0>@3 N_NET14_MMP22<0>@3_d N_VIN2_MMP22<0>@3_g N_VTAILP_MMP22<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<0>@2 N_NET13_MMP21<0>@3_d N_VIN1_MMP21<0>@2_g N_VTAILP_MMP21<0>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<0>@2 N_NET14_MMP22<0>@3_d N_VIN2_MMP22<0>@2_g N_VTAILP_MMP22<0>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<0> N_NET14_MMP22<0>_d N_VIN2_MMP22<0>_g N_VTAILP_MMP22<0>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<0> N_NET13_MMP21<0>_d N_VIN1_MMP21<0>_g N_VTAILP_MMP21<0>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP22<3>@10 N_NET14_MMP22<0>_d N_VIN2_MMP22<3>@10_g N_VTAILP_MMP22<3>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@10 N_NET13_MMP21<0>_d N_VIN1_MMP21<3>@10_g N_VTAILP_MMP21<3>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@9 N_NET14_MMP22<3>@9_d N_VIN2_MMP22<3>@9_g N_VTAILP_MMP22<3>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@9 N_NET13_MMP21<3>@9_d N_VIN1_MMP21<3>@9_g N_VTAILP_MMP21<3>@10_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@8 N_NET14_MMP22<3>@9_d N_VIN2_MMP22<3>@8_g N_VTAILP_MMP22<3>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@8 N_NET13_MMP21<3>@9_d N_VIN1_MMP21<3>@8_g N_VTAILP_MMP21<3>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@7 N_NET14_MMP22<3>@7_d N_VIN2_MMP22<3>@7_g N_VTAILP_MMP22<3>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@7 N_NET13_MMP21<3>@7_d N_VIN1_MMP21<3>@7_g N_VTAILP_MMP21<3>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@6 N_NET14_MMP22<3>@7_d N_VIN2_MMP22<3>@6_g N_VTAILP_MMP22<3>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@6 N_NET13_MMP21<3>@7_d N_VIN1_MMP21<3>@6_g N_VTAILP_MMP21<3>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@5 N_NET14_MMP22<3>@5_d N_VIN2_MMP22<3>@5_g N_VTAILP_MMP22<3>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@5 N_NET13_MMP21<3>@5_d N_VIN1_MMP21<3>@5_g N_VTAILP_MMP21<3>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@4 N_NET14_MMP22<3>@5_d N_VIN2_MMP22<3>@4_g N_VTAILP_MMP22<3>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@4 N_NET13_MMP21<3>@5_d N_VIN1_MMP21<3>@4_g N_VTAILP_MMP21<3>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@3 N_NET14_MMP22<3>@3_d N_VIN2_MMP22<3>@3_g N_VTAILP_MMP22<3>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP21<3>@3 N_NET13_MMP21<3>@3_d N_VIN1_MMP21<3>@3_g N_VTAILP_MMP21<3>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP22<3>@2 N_NET14_MMP22<3>@3_d N_VIN2_MMP22<3>@2_g N_VTAILP_MMP22<3>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP21<3>@2 N_NET13_MMP21<3>@3_d N_VIN1_MMP21<3>@2_g N_VTAILP_MMP21<3>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP16 N_NET4_MMP16_d N_NET3_MMP16_g N_VDD_MMP16_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05 NRD=0.044
+ NRS=0.026 M=1 NF=1 PAR=1
XMMP17 N_NET5_MMP17_d N_NET3_MMP17_g N_VDD_MMP17_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=3e-06 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05 NRD=0.044
+ NRS=0.026 M=1 NF=1 PAR=1
XMMP16@10 N_NET4_MMP16@10_d N_NET3_MMP16@10_g N_VDD_MMP16_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@10 N_NET5_MMP17@10_d N_NET3_MMP17@10_g N_VDD_MMP17_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@9 N_NET4_MMP16@10_d N_NET3_MMP16@9_g N_VDD_MMP16@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@9 N_NET5_MMP17@10_d N_NET3_MMP17@9_g N_VDD_MMP17@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@8 N_NET4_MMP16@8_d N_NET3_MMP16@8_g N_VDD_MMP16@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@8 N_NET5_MMP17@8_d N_NET3_MMP17@8_g N_VDD_MMP17@9_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@7 N_NET4_MMP16@8_d N_NET3_MMP16@7_g N_VDD_MMP16@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@7 N_NET5_MMP17@8_d N_NET3_MMP17@7_g N_VDD_MMP17@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@6 N_NET5_MMP17@6_d N_NET3_MMP17@6_g N_VDD_MMP16@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@6 N_NET4_MMP16@6_d N_NET3_MMP16@6_g N_VDD_MMP17@7_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@5 N_NET5_MMP17@6_d N_NET3_MMP17@5_g N_VDD_MMP17@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@5 N_NET4_MMP16@6_d N_NET3_MMP16@5_g N_VDD_MMP16@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@4 N_NET5_MMP17@4_d N_NET3_MMP17@4_g N_VDD_MMP17@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@4 N_NET4_MMP16@4_d N_NET3_MMP16@4_g N_VDD_MMP16@5_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@3 N_NET5_MMP17@4_d N_NET3_MMP17@3_g N_VDD_MMP17@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@3 N_NET4_MMP16@4_d N_NET3_MMP16@3_g N_VDD_MMP16@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP17@2 N_NET5_MMP17@2_d N_NET3_MMP17@2_g N_VDD_MMP17@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP16@2 N_NET4_MMP16@2_d N_NET3_MMP16@2_g N_VDD_MMP16@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP19 N_NET3_MMP19_d N_VBIASP_MMP19_g N_NET5_MMP17@2_d N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP18 N_NET1_MMP18_d N_VBIASP_MMP18_g N_NET4_MMP16@2_d N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP19@4 N_NET3_MMP19_d N_VBIASP_MMP19@4_g N_NET5_MMP19@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP18@4 N_NET1_MMP18_d N_VBIASP_MMP18@4_g N_NET4_MMP18@4_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP18@3 N_NET1_MMP18@3_d N_VBIASP_MMP18@3_g N_NET4_MMP18@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP19@3 N_NET3_MMP19@3_d N_VBIASP_MMP19@3_g N_NET5_MMP19@3_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP18@2 N_NET1_MMP18@3_d N_VBIASP_MMP18@2_g N_NET4_MMP18@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP19@2 N_NET3_MMP19@3_d N_VBIASP_MMP19@2_g N_NET5_MMP19@2_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-06 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP20 N_NET6_MMP20_d N_IABP_MMP20_g N_NET1_MMP20_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=1e-06 W=1e-05 AD=4.4e-12 AS=4.4e-12 PD=2.088e-05 PS=2.088e-05 NRD=0.044
+ NRS=0.044 M=1 NF=1 PAR=1
XMMP15 N_NET2_MMP15_d N_IABP_MMP15_g N_NET3_MMP15_s N_VDD_MMP14<1>_b PMOS_3P3
+ L=1e-06 W=1e-05 AD=4.4e-12 AS=4.4e-12 PD=2.088e-05 PS=2.088e-05 NRD=0.044
+ NRS=0.044 M=1 NF=1 PAR=1
XMMP3 N_VOUT_T_MMP3_d N_VSS_MMP3_g N_VOUT_MMP3_s N_VDD_MMP3_b PMOS_3P3 L=2.8e-07
+ W=2e-06 AD=8.8e-13 AS=5.2e-13 PD=4.88e-06 PS=2.52e-06 NRD=0.22 NRS=0.13 M=1
+ NF=1 PAR=1
XMMP3@12 N_VOUT_T_MMP3@12_d N_VSS_MMP3@12_g N_VOUT_MMP3_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@11 N_VOUT_T_MMP3@12_d N_VSS_MMP3@11_g N_VOUT_MMP3@11_s N_VDD_MMP3_b
+ PMOS_3P3 L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMP3@10 N_VOUT_T_MMP3@10_d N_VSS_MMP3@10_g N_VOUT_MMP3@11_s N_VDD_MMP3_b
+ PMOS_3P3 L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06
+ NRD=0.13 NRS=0.13 M=1 NF=1 PAR=1
XMMP3@9 N_VOUT_T_MMP3@10_d N_VSS_MMP3@9_g N_VOUT_MMP3@9_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@8 N_VOUT_T_MMP3@8_d N_VSS_MMP3@8_g N_VOUT_MMP3@9_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@7 N_VOUT_T_MMP3@8_d N_VSS_MMP3@7_g N_VOUT_MMP3@7_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@6 N_VOUT_T_MMP3@6_d N_VSS_MMP3@6_g N_VOUT_MMP3@7_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@5 N_VOUT_T_MMP3@6_d N_VSS_MMP3@5_g N_VOUT_MMP3@5_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@4 N_VOUT_T_MMP3@4_d N_VSS_MMP3@4_g N_VOUT_MMP3@5_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@3 N_VOUT_T_MMP3@4_d N_VSS_MMP3@3_g N_VOUT_MMP3@3_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=5.2e-13 AS=5.2e-13 PD=2.52e-06 PS=2.52e-06 NRD=0.13
+ NRS=0.13 M=1 NF=1 PAR=1
XMMP3@2 N_VOUT_T_MMP3@2_d N_VSS_MMP3@2_g N_VOUT_MMP3@3_s N_VDD_MMP3_b PMOS_3P3
+ L=2.8e-07 W=2e-06 AD=8.8e-13 AS=5.2e-13 PD=4.88e-06 PS=2.52e-06 NRD=0.22
+ NRS=0.13 M=1 NF=1 PAR=1
D432_noxref N_VSS_MMN25<4>_b N_VDD_D432_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D433_noxref N_VSS_MMN25<4>_b N_VDD_D433_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D434_noxref N_VSS_MMN25<4>_b N_VDD_D434_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D435_noxref N_VSS_MMN25<4>_b N_VDD_D435_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D436_noxref N_VSS_MMN25<4>_b N_VDD_D436_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D437_noxref N_VSS_MMN25<4>_b N_VDD_D437_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D438_noxref N_VSS_MMN25<4>_b N_VDD_D438_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D439_noxref N_VSS_MMN25<4>_b N_VDD_D439_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D440_noxref N_VSS_MMN25<4>_b N_VDD_D440_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D441_noxref N_VSS_MMN25<4>_b N_VDD_D441_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D442_noxref N_VSS_MMN25<4>_b N_VDD_D442_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D443_noxref N_VSS_MMN25<4>_b N_VDD_D443_noxref_neg np_3p3  AREA=2.5392e-11
+ PJ=0.0001058 M=1
D444_noxref N_VSS_MMN25<4>_b N_noxref_5005_D444_noxref_neg np_3p3 
+ AREA=2.5392e-11 PJ=0.0001058 M=1
D445_noxref N_VSS_MMN25<4>_b N_noxref_5005_D445_noxref_neg np_3p3 
+ AREA=2.5392e-11 PJ=0.0001058 M=1
D446_noxref N_VSS_MMN25<4>_b N_VDD_D446_noxref_neg np_3p3  AREA=1.896e-11
+ PJ=7.9e-05 M=1
D447_noxref N_VSS_MMN25<4>_b N_VDD_D447_noxref_neg np_3p3  AREA=1.896e-11
+ PJ=7.9e-05 M=1
D448_noxref N_VSS_MMN25<4>_b N_VDD_D448_noxref_neg np_3p3  AREA=2.01408e-11
+ PJ=8.392e-05 M=1
D449_noxref N_VSS_MMN25<4>_b N_VDD_D449_noxref_neg np_3p3  AREA=2.028e-11
+ PJ=8.45e-05 M=1
D450_noxref N_VSS_MMN25<4>_b N_VDD_D450_noxref_neg np_3p3  AREA=2.1055e-11
+ PJ=8.54e-05 M=1
D451_noxref N_VSS_MMN25<4>_b N_VDD_D451_noxref_neg np_3p3  AREA=2.02944e-11
+ PJ=8.456e-05 M=1
D452_noxref N_VSS_MMN25<4>_b N_VDD_D452_noxref_neg np_3p3  AREA=2.54111e-10
+ PJ=0.00025344 M=1
D453_noxref N_VSS_MMN25<4>_b N_VDD_MMP14<1>_b nwp_3p3  AREA=4.95832e-09
+ PJ=0.00042095 M=1
D454_noxref N_VSS_MMN25<4>_b N_VDD_MMP3_b nwp_3p3  AREA=3.04006e-10 PJ=8.324e-05
+ M=1
XCC4 N_NET1_CC4_pos N_VOUT_CC4_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05 M=1
XCC4__2 N_NET1_CC4__2_pos N_VOUT_CC4__2_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05
+ M=1
XCC5 N_NET6_CC5_pos N_VOUT_CC5_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05 M=1
XCC5__2 N_NET6_CC5__2_pos N_VOUT_CC5__2_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05
+ M=1
XCC4__3 N_NET1_CC4__3_pos N_VOUT_CC4__3_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05
+ M=1
XCC5__3 N_NET6_CC5__3_pos N_VOUT_CC5__3_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05
+ M=1
XCC5__4 N_NET6_CC5__4_pos N_VOUT_CC5__4_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05
+ M=1
XCC4__4 N_NET1_CC4__4_pos N_VOUT_CC4__4_neg mim_2p0fF  PAR=1 L=2.5e-05 W=2.5e-05
+ M=1
XMMP14<1> N_VOUT_MMP14<1>_d N_NET1_MMP14<1>_g N_VDD_MMP14<1>_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05 PS=1.052e-05
+ NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@7 N_VOUT_MMP14<0>@7_d N_NET1_MMP14<0>@7_g N_VDD_MMP14<1>_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@6 N_VOUT_MMP14<0>@7_d N_NET1_MMP14<0>@6_g N_VDD_MMP14<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@5 N_VOUT_MMP14<0>@5_d N_NET1_MMP14<0>@5_g N_VDD_MMP14<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@4 N_VOUT_MMP14<0>@5_d N_NET1_MMP14<0>@4_g N_VDD_MMP14<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@3 N_VOUT_MMP14<0>@3_d N_NET1_MMP14<0>@3_g N_VDD_MMP14<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@2 N_VOUT_MMP14<0>@3_d N_NET1_MMP14<0>@2_g N_VDD_MMP14<0>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0> N_VOUT_MMP14<0>_d N_NET1_MMP14<0>_g N_VDD_MMP14<0>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<0>@8 N_VOUT_MMP14<0>_d N_NET1_MMP14<0>@8_g N_VDD_MMP14<0>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<1>@7 N_VOUT_MMP14<1>@7_d N_NET1_MMP14<1>@7_g N_VDD_MMP14<0>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<1>@6 N_VOUT_MMP14<1>@7_d N_NET1_MMP14<1>@6_g N_VDD_MMP14<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<1>@5 N_VOUT_MMP14<1>@5_d N_NET1_MMP14<1>@5_g N_VDD_MMP14<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<1>@4 N_VOUT_MMP14<1>@5_d N_NET1_MMP14<1>@4_g N_VDD_MMP14<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<1>@3 N_VOUT_MMP14<1>@3_d N_NET1_MMP14<1>@3_g N_VDD_MMP14<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP14<1>@2 N_VOUT_MMP14<1>@3_d N_NET1_MMP14<1>@2_g N_VDD_MMP14<1>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP13<2> N_VDD_MMP13<2>_d N_VDD_MMP13<2>_g N_VDD_MMP13<2>_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05 PS=2.088e-05
+ NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP13<1>@5 N_VDD_MMP13<1>@5_d N_VDD_MMP13<1>@5_g N_VDD_MMP13<2>_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1>@4 N_VDD_MMP13<1>@4_d N_VDD_MMP13<1>@4_g N_VDD_MMP13<1>@5_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1>@3 N_VDD_MMP13<1>@3_d N_VDD_MMP13<1>@3_g N_VDD_MMP13<1>@4_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1>@2 N_VDD_MMP13<1>@2_d N_VDD_MMP13<1>@2_g N_VDD_MMP13<1>@3_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1> N_VDD_MMP13<1>_d N_VDD_MMP13<1>_g N_VDD_MMP13<1>@2_d N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1>@8 N_VDD_MMP13<1>@8_d N_VDD_MMP13<1>@8_g N_VDD_MMP13<1>_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1>@7 N_VDD_MMP13<1>@7_d N_VDD_MMP13<1>@7_g N_VDD_MMP13<1>@8_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<1>@6 N_VDD_MMP13<1>@6_d N_VDD_MMP13<1>@6_g N_VDD_MMP13<1>@7_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0>@5 N_VDD_MMP13<0>@5_d N_VDD_MMP13<0>@5_g N_VDD_MMP13<1>@6_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0>@4 N_VDD_MMP13<0>@4_d N_VDD_MMP13<0>@4_g N_VDD_MMP13<0>@5_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0>@3 N_VDD_MMP13<0>@3_d N_VDD_MMP13<0>@3_g N_VDD_MMP13<0>@4_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0>@2 N_VDD_MMP13<0>@2_d N_VDD_MMP13<0>@2_g N_VDD_MMP13<0>@3_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0> N_VDD_MMP13<0>_d N_VDD_MMP13<0>_g N_VDD_MMP13<0>@2_d N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0>@8 N_VDD_MMP13<0>@8_d N_VDD_MMP13<0>@8_g N_VDD_MMP13<0>_d
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<0>@7 N_VDD_MMP13<0>@7_d N_VDD_MMP13<0>@7_g N_VDD_MMP13<0>@7_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMP13<0>@6 N_VDD_MMP13<0>@7_s N_VDD_MMP13<0>@6_g N_VDD_MMP13<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@5 N_VDD_MMP13<0>@6_s N_VDD_MMN26<2>@5_g N_VDD_MMN26<2>@5_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@4 N_VDD_MMN26<2>@5_s N_VDD_MMN26<2>@4_g N_VDD_MMN26<2>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@3 N_VDD_MMN26<2>@4_s N_VDD_MMN26<2>@3_g N_VDD_MMN26<2>@3_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@2 N_VDD_MMN26<2>@3_s N_VDD_MMN26<2>@2_g N_VDD_MMN26<2>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2> N_VDD_MMN26<2>@2_s N_VDD_MMN26<2>_g N_VDD_MMN26<2>_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@8 N_VDD_MMN26<2>_s N_VDD_MMN26<2>@8_g N_VDD_MMN26<2>@8_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@7 N_VDD_MMN26<2>@8_s N_VDD_MMN26<2>@7_g N_VDD_MMN26<2>@7_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<2>@6 N_VDD_MMN26<2>@7_s N_VDD_MMN26<2>@6_g N_VDD_MMN26<2>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<1>@7 N_VDD_MMN26<2>@6_s N_VDD_MMN26<1>@7_g N_VDD_MMN26<1>@7_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<1>@6 N_VDD_MMN26<1>@7_s N_VDD_MMN26<1>@6_g N_VDD_MMN26<1>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<1>@5 N_VDD_MMN26<1>@6_s N_VDD_MMN26<1>@5_g N_VDD_MMN26<1>@5_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<1>@4 N_VDD_MMN26<1>@5_s N_VDD_MMN26<1>@4_g N_VDD_MMN26<1>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<1>@3 N_VDD_MMN26<1>@4_s N_VDD_MMN26<1>@3_g N_VDD_MMN26<1>@3_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<1>@2 N_VDD_MMN26<1>@2_d N_VDD_MMN26<1>@2_g N_VDD_MMN26<1>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=4.4e-12 PD=1.052e-05
+ PS=2.088e-05 NRD=0.026 NRS=0.044 M=1 NF=1 PAR=1
XMMN26<1> N_VDD_MMN26<1>@2_s N_VDD_MMN26<1>_g N_VDD_MMN26<1>_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0>@7 N_VDD_MMN26<1>_s N_VDD_MMN26<0>@7_g N_VDD_MMN26<0>@7_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0>@6 N_VDD_MMN26<0>@7_s N_VDD_MMN26<0>@6_g N_VDD_MMN26<0>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0>@5 N_VDD_MMN26<0>@6_s N_VDD_MMN26<0>@5_g N_VDD_MMN26<0>@5_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0>@4 N_VDD_MMN26<0>@5_s N_VDD_MMN26<0>@4_g N_VDD_MMN26<0>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0>@3 N_VDD_MMN26<0>@4_s N_VDD_MMN26<0>@3_g N_VDD_MMN26<0>@3_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0>@2 N_VDD_MMN26<0>@3_s N_VDD_MMN26<0>@2_g N_VDD_MMN26<0>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMN26<0> N_VDD_MMN26<0>@2_s N_VDD_MMN26<0>_g N_VDD_MMN26<0>_s N_VDD_MMP14<1>_b
+ PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05 PS=1.052e-05
+ NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<2>@7 N_VDD_MMN26<0>_s N_VDD_MMP13<2>@7_g N_VDD_MMP13<2>@7_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<2>@6 N_VDD_MMP13<2>@7_s N_VDD_MMP13<2>@6_g N_VDD_MMP13<2>@6_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<2>@5 N_VDD_MMP13<2>@6_s N_VDD_MMP13<2>@5_g N_VDD_MMP13<2>@5_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<2>@4 N_VDD_MMP13<2>@5_s N_VDD_MMP13<2>@4_g N_VDD_MMP13<2>@4_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<2>@3 N_VDD_MMP13<2>@4_s N_VDD_MMP13<2>@3_g N_VDD_MMP13<2>@3_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=2.6e-12 AS=2.6e-12 PD=1.052e-05
+ PS=1.052e-05 NRD=0.026 NRS=0.026 M=1 NF=1 PAR=1
XMMP13<2>@2 N_VDD_MMP13<2>@3_s N_VDD_MMP13<2>@2_g N_VDD_MMP13<2>@2_s
+ N_VDD_MMP14<1>_b PMOS_3P3 L=3e-07 W=1e-05 AD=4.4e-12 AS=2.6e-12 PD=2.088e-05
+ PS=1.052e-05 NRD=0.044 NRS=0.026 M=1 NF=1 PAR=1
*
.include "opamp2_hspice.pex.netlist.OPAMP2_NODW.pxi"
*
.ends
*
*
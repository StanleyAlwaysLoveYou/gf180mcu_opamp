.include /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/stanleylin/silicon-env/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical


.param  sw_stat_mismatch = 0
.param  sw_stat_global = 0

.include ../netlist/Programmable_2stage_opamp_wo_res_pex.spice
X1 vout vout_t vbiasp vbiasn vin2 vin1 vprog vss vdd opamp2

V1 vdd GND 3.3
V2 vss GND 0
V3 vin1 GND dc 0.8 ac 1
V4 vin2 GND dc 0.8 ac 0 
V5 vprog GND dc 0
V6 vbiasp GND dc 0.9
V7 vbiasn GND dc 1



.save i(v1)
.save i(v2)
.save i(v3)
.save i(v4)
.save i(v5)
.save all

.control

let begin = 1
let step = 0.1
let final = 1
let test = begin
let cnt = 0

set color0 = white
set color1 = black
set hcopydevtype = svg
setcs svg_stropts = ( black Arial Arial )

set nolegend

set gain = ' '
set phasedeg = ' '
let ind = ((final-begin)/step)
let dc_gains = vector(ind)
let bandwidths = vector(ind)
let phase_margins = vector(ind)
let power = vector(ind)


let test = begin
while test le final

    alter @v5[dc] = test
    print @v5[dc]
    let test = test + step

    op

    let ic = v1#branch
    let power[cnt] = 3.3*(-ic)
    print power[cnt]
    let cnt = cnt + 1

end




let test = begin
let cnt = 0

while test le final

    alter @v5[dc] = test
    print @v5[dc]
    let test = test + step

    ac dec 10 1 300MEG

    let phase = {57.29*vp(vout)}-180
    set gain = ( $gain db({$curplot}.vout) )
    set phasedeg = ( $phasedeg ({$curplot}.phase) )
    let dbvout = db(vout)


    meas ac dc_gain find dbvout at=10
    meas ac bandwidth when dbvout=0
    let pm = phase +180
    meas ac phase_margin find pm at=bandwidth

    let dc_gains[cnt] = dc_gain
    let bandwidths[cnt] = bandwidth
    let phase_margins[cnt] = phase_margin

    let cnt = cnt + 1
    

end



plot $gain xlabel Frequency(Hz) ylabel Gain(db) title Gain(dB)
plot $phasedeg xlabel Frequency(Hz) ylabel Phase(deg) title Phase(deg)
plot dc_gains vs power xlabel Power(mW) ylabel Gain(db) title OTA_2stage_Gain_vs_Power
plot bandwidths vs power xlabel Power(mW) ylabel Frequency(Hz) title OTA_2stage_GBW_vs_Power
plot phase_margins vs power xlabel Power(mW) ylabel Phase_margin title OTA_2stage_PM_vs_Power


hardcopy ../output/Gain.svg $gain xlabel Frequency(Hz) ylabel Gain(db) title 'OTA_2stage Gain'
hardcopy ../output/Phase.svg $phasedeg xlabel Frequency(Hz) ylabel Phase(deg) title 'OTA_2stage Phase'
hardcopy ../output/Gain_vs_Power.svg dc_gains vs power xlabel Power(mW) ylabel Gain(db) title 'OTA_2stage_Gain_vs_Power'
hardcopy ../output/GBW_vs_Power.svg bandwidths vs power xlabel Power(mW) ylabel Frequency(Hz) title 'OTA_2stage_GBW_vs_Power'
hardcopy ../output/PM_vs_Power.svg phase_margins vs power xlabel Power(mW) ylabel Phase_margin title 'OTA_2stage_PM_vs_Power'

print power

.endc


.GLOBAL GND

.end
